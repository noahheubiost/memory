-- # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # #
-- #                                                                     #
-- #      Hardware description by Lukas Leuenberger l1leuenb@hsr.ch      #
-- #                                                                     #
-- #                            Created: 12.12.2019                      #
-- #                        Last modified: 12.12.2019                     #
-- #                                                                     #
-- #          Copyright by Hochschule fuer Technik in Rapperswil         #
-- #                                                                     #
-- #                                                                     #
-- # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # #

------------------------------------------------------------------------------------------------
-- Library declarations
------------------------------------------------------------------------------------------------
-- Standard library ieee	
library ieee;
-- This package defines the basic std_logic data types and a few functions.								
use ieee.std_logic_1164.all;
-- This package provides arithmetic functions for vectors.		
use ieee.numeric_std.all;
-- This package provides functions for the calcualtion with real values.
use ieee.math_real.all;
-- This package provides file specific functions.
use std.textio.all;
-- This package provides file specific functions for the std_logic types.
use ieee.std_logic_textio.all;

------------------------------------------------------------------------------------------------
-- Entity declarations
------------------------------------------------------------------------------------------------
entity bmpImage is
	generic(
		imSizeH_g : integer := 256; --output picture size
		imSizeV_g : integer := 256; --output picture size
		-- bus size
		rowSize_g      : integer := 8;
		colSize_g      : integer := 8
	);
	port(
		-- Reset und Clock
		resetn     : in  std_logic;     -- Synchronous Negative Reset
		clk        : in  std_logic;     -- Clock
		-- FPGA Image out
		row_out    : out unsigned(rowSize_g - 1 downto 0);
		col_out    : out unsigned(colSize_g - 1 downto 0);
		d_out      : out std_logic_vector(15 downto 0);
		strobe_out : out std_logic
	);
end entity bmpImage;

---------------------------------------------------------------------
-- Architecture declarations
---------------------------------------------------------------------
architecture RTL of bmpImage is	
	------------------------------------------------------------------------------------------------
	-- internal types
	------------------------------------------------------------------------------------------------
	type rom_type is array (0 to (imSizeH_g * imSizeV_g) - 1) of std_logic_vector(15 downto 0);	
	
	------------------------------------------------------------------------------------------------
	-- Internal constants
	------------------------------------------------------------------------------------------------
	constant blockrom : rom_type := (x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFFF",x"FFFF",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",
									 x"FFDF",x"FFDF",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",
									 x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",
									 x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"FFDF",x"F7DF",
									 x"F7DF",x"F7DF",x"F7BF",x"F7BF",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F79E",x"F79E",
									 x"F79E",x"F79E",x"EF7D",x"EF7D",x"EF7E",x"EF7E",x"EF7E",x"EF7E",x"EF7E",x"EF7D",
									 x"EF7D",x"EF7E",x"EF7E",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",
									 x"EF7D",x"EF9D",x"EF9D",x"EF9E",x"EF9E",x"F79E",x"F7BE",x"F79E",x"F7BE",x"FFBE",
									 x"FFDF",x"FFDF",x"FFDF",x"FFFF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDF",
									 x"FFDF",x"FFDE",x"FFDE",x"F7BE",x"F7BE",x"F7BE",x"F79E",x"F79E",x"F79E",x"EF9E",
									 x"EF7E",x"EF7E",x"EF7D",x"EF7D",x"EF5D",x"EF5D",x"E75C",x"E75C",x"E75C",x"E75C",
									 x"E75C",x"EF5C",x"EF3C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",
									 x"E73C",x"E73C",x"E71B",x"E71B",x"EF1B",x"E71B",x"E73B",x"E73C",x"E73B",x"E73C",
									 x"E73D",x"EF5D",x"EF5D",x"EF7D",x"EF7D",x"F79D",x"F79E",x"F79E",x"F7BE",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDE",x"FFDE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDF",x"FFDF",x"FFDF",x"FFBE",x"F7BF",x"FFBE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",
									 x"F77D",x"F75C",x"F73B",x"F71A",x"F6D9",x"EED9",x"EEB8",x"EE97",x"EE97",x"EE76",
									 x"EE56",x"EE35",x"EE34",x"EE34",x"EE34",x"EE33",x"EE13",x"EE13",x"EE13",x"EE12",
									 x"EE12",x"EE12",x"EE12",x"EE13",x"EE13",x"EE13",x"E614",x"E614",x"E615",x"E635",
									 x"E635",x"E655",x"E656",x"E677",x"E678",x"E699",x"E6B9",x"EEDA",x"E6FB",x"E73C",
									 x"E75D",x"E75D",x"EF7C",x"EF7D",x"EF7D",x"F79D",x"F79D",x"F7BE",x"F7BF",x"F7DF",
									 x"F7DF",x"F7DF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F7FF",x"F7DF",x"F7DF",x"F7DF",x"F7BF",x"F79E",
									 x"F77D",x"EF5D",x"EF5C",x"EF3C",x"EF5C",x"F71A",x"F6D9",x"EE97",x"EE55",x"EDF3",
									 x"EDB1",x"ED6F",x"F52D",x"ECEC",x"E4CA",x"ECA9",x"EC88",x"EC68",x"EC67",x"EC67",
									 x"EC46",x"EC25",x"EC24",x"EC24",x"EC24",x"EC04",x"EC04",x"EC24",x"EC24",x"EC24",
									 x"EC45",x"EC66",x"EC67",x"EC68",x"EC88",x"E489",x"DCAA",x"E4EB",x"E50D",x"E52E",
									 x"E570",x"EDB2",x"E5D3",x"E614",x"E656",x"E698",x"E6B9",x"DEDA",x"E6DB",x"DEDB",
									 x"DEFB",x"E71C",x"E73D",x"E73D",x"EF5E",x"EF7E",x"EF7E",x"EF9E",x"F7BE",x"F7DE",
									 x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"F7BF",
									 x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F77D",x"F75C",x"F71B",x"EED9",x"EE97",x"EE56",
									 x"E635",x"EDF2",x"EDB0",x"ED6F",x"E50D",x"E4EB",x"ECCA",x"ECA9",x"ECA8",x"EC67",
									 x"EC46",x"EC45",x"EC45",x"EC24",x"F424",x"F423",x"F423",x"F422",x"F422",x"F402",
									 x"F402",x"F402",x"F402",x"F401",x"F401",x"F402",x"F422",x"F423",x"EC23",x"EC24",
									 x"EC45",x"EC45",x"EC45",x"EC66",x"EC87",x"EC88",x"ECA9",x"ECCA",x"E4EC",x"E50D",
									 x"E54E",x"DD70",x"E5B2",x"E5F4",x"DE16",x"DE37",x"DE78",x"E6DA",x"E6FB",x"E71C",
									 x"E71B",x"E71B",x"E71C",x"E73C",x"E75D",x"EF7D",x"F79E",x"F79E",x"F7BE",x"F7BE",
									 x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDF",x"F7BE",x"F7BE",x"F7BD",x"F77C",x"F75B",x"F73A",x"F71A",
									 x"F6D8",x"F676",x"F655",x"F5F2",x"ED90",x"ED4E",x"ED0D",x"ECEA",x"ECC9",x"ECA8",
									 x"EC87",x"EC66",x"EC66",x"EC45",x"EC45",x"EC45",x"EC44",x"EC44",x"EC44",x"F444",
									 x"F444",x"F444",x"F443",x"F443",x"F463",x"F443",x"F443",x"F443",x"F443",x"F443",
									 x"F443",x"F463",x"F463",x"F463",x"F463",x"F464",x"F464",x"F464",x"F443",x"EC44",
									 x"EC44",x"EC45",x"EC65",x"EC86",x"EC86",x"EC87",x"ECA9",x"E4CA",x"E4EB",x"ED2D",
									 x"E54E",x"ED90",x"E5D1",x"E634",x"E655",x"E676",x"E6B8",x"E6B8",x"DEB9",x"DEDA",
									 x"DEFC",x"E71D",x"E75D",x"EF5D",x"EF7D",x"EF7D",x"F79E",x"F7BE",x"F7BE",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDE",x"FFBE",x"FFBE",x"FFBE",x"FFBE",
									 x"F79D",x"FF5B",x"F6F8",x"F696",x"F633",x"EDD1",x"E56F",x"ED0D",x"ECCB",x"ECA9",
									 x"EC67",x"EC66",x"F466",x"EC45",x"EC44",x"EC44",x"EC44",x"F464",x"F464",x"F463",
									 x"F463",x"F463",x"F463",x"F462",x"F462",x"F463",x"F463",x"F483",x"F483",x"F483",
									 x"F483",x"F483",x"F483",x"F483",x"F483",x"F483",x"F483",x"F483",x"F4A3",x"F483",
									 x"F483",x"F482",x"F482",x"F483",x"F483",x"F483",x"F483",x"F483",x"F463",x"F463",
									 x"F464",x"EC44",x"EC44",x"EC65",x"EC45",x"EC66",x"EC87",x"ECA8",x"E4C9",x"E4EB",
									 x"E52C",x"E56E",x"DDB1",x"E5F3",x"E635",x"E678",x"E6BA",x"E6FB",x"E6FA",x"E6FB",
									 x"E71B",x"E71C",x"E73D",x"EF5D",x"F79D",x"F7BE",x"F7DF",x"FFFF",x"FFDF",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F7DE",x"F7BE",
									 x"F7BF",x"F7BD",x"F77C",x"F71A",x"F6D9",x"F697",x"EE55",x"EE12",x"EDB0",x"ED2D",
									 x"ECEB",x"ECA9",x"E487",x"EC46",x"EC25",x"EC24",x"EC23",x"EC23",x"F422",x"F443",
									 x"F442",x"F442",x"F462",x"F462",x"F483",x"F483",x"F4A3",x"F4C3",x"F4C3",x"F4C3",
									 x"F4C3",x"F4C3",x"F4C3",x"F4C3",x"F4C3",x"F4C3",x"F4C3",x"F4C3",x"F4C3",x"F4C3",
									 x"F4E3",x"FCE4",x"F4C3",x"F4C3",x"F4C4",x"F4C3",x"F4C3",x"F4C3",x"F4C3",x"F4C3",
									 x"F4C3",x"F4A3",x"FCA3",x"FCA3",x"F4A3",x"F483",x"F483",x"F483",x"F463",x"F463",
									 x"F463",x"F463",x"F443",x"F444",x"EC44",x"EC65",x"E466",x"EC87",x"E4A9",x"E4CB",
									 x"E50D",x"DD70",x"DDB3",x"DDF4",x"DE15",x"DE36",x"DE98",x"DEBA",x"DEFC",x"E71C",
									 x"DF3C",x"E73C",x"E77D",x"EF9E",x"F79E",x"FFBE",x"F7DF",x"F7DF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFDF",x"F7DF",x"F7DF",x"F7BE",x"F77D",x"F75C",x"F75B",x"F6D8",x"EE55",
									 x"F5D1",x"F56E",x"ED0B",x"ECA9",x"EC88",x"EC66",x"EC45",x"EC44",x"F423",x"EC44",
									 x"F444",x"F463",x"F463",x"F463",x"F483",x"F483",x"F483",x"FCA3",x"F4A3",x"F4A3",
									 x"F4C3",x"F4C3",x"F4E4",x"F4E4",x"FCE4",x"FCE4",x"FCE3",x"FCE4",x"FCE4",x"FCE4",
									 x"FD04",x"FD04",x"FD04",x"FD04",x"FD04",x"FD04",x"FD04",x"FD04",x"FCE4",x"F4E4",
									 x"F4E4",x"FCE4",x"FCE3",x"F4E3",x"F4E3",x"F4E3",x"FCE3",x"FCE3",x"FCE3",x"FCC3",
									 x"F4C3",x"F4A3",x"F4A3",x"F4A3",x"FCA3",x"F4A3",x"F483",x"F483",x"F483",x"F483",
									 x"F463",x"EC63",x"EC63",x"EC64",x"F444",x"EC65",x"EC67",x"E4A9",x"E4CA",x"E50C",
									 x"DD2E",x"DD91",x"E614",x"E677",x"DE98",x"DEBA",x"DEDB",x"DEDB",x"DF1C",x"DF3D",
									 x"E75D",x"EF9E",x"F7BE",x"F7BF",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"FFDF",x"FFDE",x"FFDE",x"FFBE",x"F79E",
									 x"F75B",x"EEB8",x"EE55",x"F5F2",x"ED6F",x"ED0C",x"F4CA",x"F487",x"F446",x"F424",
									 x"F423",x"F422",x"F442",x"FC42",x"F442",x"F462",x"F482",x"FCA2",x"F4A2",x"F4A3",
									 x"F4C4",x"FCC4",x"FCC4",x"FCE4",x"F4E3",x"F4E3",x"F504",x"F504",x"F504",x"FD24",
									 x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",
									 x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD23",
									 x"FD23",x"FD23",x"FD23",x"FD03",x"FD03",x"FD03",x"FD03",x"FCE3",x"FCE3",x"F4E3",
									 x"F4E3",x"F4C3",x"F4C3",x"F4A3",x"F4A3",x"F4A3",x"FCA3",x"F4A3",x"F483",x"F462",
									 x"FC42",x"F442",x"F443",x"EC44",x"EC45",x"E465",x"EC87",x"ECC9",x"E50C",x"E54E",
									 x"DD91",x"E5F3",x"DE16",x"DE58",x"E6DA",x"DEFB",x"DF1B",x"DF3C",x"E73C",x"EF5D",
									 x"F77D",x"F79E",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDE",x"FFDF",x"FFDF",
									 x"FFBE",x"FF9D",x"FF7B",x"FF19",x"F6D8",x"F696",x"F613",x"ED6F",x"ED0C",x"F488",
									 x"EC26",x"EC05",x"EC04",x"EC03",x"EC03",x"F443",x"F463",x"F483",x"F482",x"F4A3",
									 x"FCA3",x"F4A2",x"F4C2",x"FCE3",x"FD03",x"FD04",x"FD04",x"FD04",x"FD04",x"FD24",
									 x"F524",x"F524",x"F524",x"FD24",x"FD24",x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",
									 x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",
									 x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",x"FD43",x"FD44",x"FD44",x"FD43",
									 x"FD23",x"FD24",x"FD23",x"FD23",x"FD23",x"FD23",x"F503",x"F503",x"FD03",x"FCE3",
									 x"FCE4",x"FCE4",x"FCC4",x"FCC4",x"FCC3",x"FCA3",x"FCA2",x"F482",x"F483",x"F483",
									 x"F483",x"EC63",x"F422",x"F443",x"EC45",x"E466",x"E4A9",x"ED0B",x"E56F",x"E591",
									 x"E614",x"DE56",x"DE77",x"DE98",x"DEBA",x"E6DA",x"E71B",x"EF5D",x"EF7E",x"F7BF",
									 x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFDF",x"F7BE",x"F7DE",x"FFBE",x"FF9E",x"FF5C",x"FF3A",x"F6D8",x"EE13",
									 x"E56F",x"ECEB",x"EC68",x"EC25",x"EC24",x"F444",x"F423",x"F443",x"F443",x"F463",
									 x"F482",x"F483",x"F4A3",x"F4C3",x"F4C3",x"F4C4",x"FCC4",x"F4E4",x"FD04",x"FD23",
									 x"FD24",x"FD24",x"FD25",x"FD45",x"FD45",x"FD44",x"FD44",x"FD64",x"FD64",x"FD64",
									 x"FD65",x"FD65",x"FD65",x"FD85",x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",
									 x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",x"FD64",x"FD64",x"FD84",x"FD84",
									 x"FD84",x"FD84",x"FD64",x"FD64",x"FD64",x"FD64",x"FD64",x"FD64",x"FD64",x"FD44",
									 x"FD64",x"FD44",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD04",x"FD03",
									 x"FCE3",x"FCE3",x"F4E3",x"F4C3",x"F4C3",x"F4C3",x"F4A2",x"F482",x"F483",x"F463",
									 x"F463",x"F443",x"EC44",x"EC65",x"E466",x"E4A8",x"DCEC",x"DD50",x"DDB3",x"DE16",
									 x"DE78",x"DE99",x"DEB9",x"DEDA",x"DEDB",x"DF1C",x"EF5D",x"F79E",x"FFDF",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F7FF",x"FFDF",x"FFDF",x"F7BF",
									 x"FF7D",x"FF1B",x"F6B7",x"F634",x"F5B1",x"ED2D",x"ECA9",x"F466",x"F424",x"F423",
									 x"F423",x"EC43",x"EC63",x"F463",x"F483",x"F4A2",x"F4C2",x"F4A3",x"F4C3",x"FD04",
									 x"F504",x"F504",x"FD04",x"F504",x"F524",x"FD44",x"FD44",x"FD44",x"FD45",x"FD65",
									 x"FD65",x"FD65",x"FD64",x"FD84",x"FD84",x"FD84",x"FD85",x"FD85",x"FD85",x"FD85",
									 x"FD85",x"FD85",x"FD85",x"FD85",x"FD85",x"FD85",x"FD85",x"FD85",x"FD85",x"FD85",
									 x"FD85",x"FD85",x"FD85",x"FD84",x"FD85",x"FD85",x"FD84",x"FD84",x"FD84",x"FD84",
									 x"FD84",x"FD84",x"FD64",x"FD84",x"FD64",x"FD64",x"FD64",x"FD64",x"FD44",x"FD44",
									 x"FD44",x"FD44",x"FD43",x"FD43",x"FD23",x"F523",x"F523",x"F523",x"F503",x"F503",
									 x"FD03",x"F4E2",x"F4C2",x"FCC2",x"F4C3",x"F4A3",x"F483",x"F483",x"F463",x"F463",
									 x"F463",x"F464",x"EC87",x"E4CA",x"E50D",x"E54F",x"DDD3",x"D615",x"D657",x"D699",
									 x"D6BB",x"D6FC",x"DF1C",x"E75D",x"EF9E",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FFDF",
									 x"FFFF",x"F7FF",x"F7DF",x"FFBE",x"FF7D",x"FF1B",x"F697",x"F613",x"E54D",x"E4A9",
									 x"EC47",x"EC25",x"EC04",x"EC23",x"F443",x"F463",x"F463",x"F483",x"F483",x"F4A3",
									 x"F4C3",x"F4E3",x"F4E3",x"FD03",x"FD04",x"FD04",x"FD04",x"FD24",x"FD44",x"FD44",
									 x"FD44",x"FD64",x"FD64",x"FD64",x"FD65",x"FD85",x"FD85",x"FD85",x"FD85",x"FD85",
									 x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",
									 x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",
									 x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FD85",x"FD85",x"FD85",x"FD85",x"FD84",x"FD84",
									 x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",x"FD64",x"FD84",x"FD84",x"FD64",x"FD64",
									 x"FD64",x"FD43",x"FD43",x"FD43",x"FD23",x"FD23",x"FD23",x"F503",x"FD03",x"F503",
									 x"F4E3",x"F4E3",x"F4C3",x"F4C3",x"F4A3",x"F4A3",x"F462",x"F463",x"EC44",x"EC45",
									 x"E466",x"E487",x"DCEB",x"DD4E",x"DDB1",x"DE15",x"DE98",x"D69A",x"CEBA",x"D6DC",
									 x"DEFC",x"EF3C",x"F77D",x"F7BE",x"F7DF",x"FFFF",x"FFFE",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F7DF",x"F7DF",x"FFDF",x"FFBE",x"FF3B",x"FED8",
									 x"F634",x"ED8F",x"ECEB",x"EC88",x"EC66",x"EC44",x"EC23",x"EC43",x"F443",x"F462",
									 x"F482",x"FCA2",x"F4C2",x"FCC3",x"FCE4",x"FCE4",x"FD04",x"FD04",x"FD24",x"FD24",
									 x"FD24",x"FD24",x"FD44",x"FD44",x"FD65",x"FD65",x"FD65",x"FD85",x"FD85",x"FD85",
									 x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",
									 x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",
									 x"FDC5",x"FDC5",x"FDC5",x"FDC6",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",
									 x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA4",x"FD84",x"FDA4",x"FDA4",
									 x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD84",x"FD64",x"FD64",x"FD64",
									 x"FD64",x"FD44",x"FD44",x"FD44",x"FD24",x"FD23",x"FD03",x"FD03",x"F503",x"F4E3",
									 x"F4E3",x"F4C3",x"FCC3",x"FCA2",x"F482",x"F483",x"EC63",x"EC63",x"EC66",x"E487",
									 x"E4A9",x"E50C",x"DD90",x"DDD3",x"D616",x"D679",x"D69A",x"DEBA",x"DEDB",x"E73C",
									 x"E77D",x"F7BF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F7FF",x"F7DF",
									 x"F7DF",x"F7BE",x"FF9E",x"FF1B",x"FE97",x"FE33",x"F58E",x"ECC7",x"EC25",x"F3E3",
									 x"F403",x"EC22",x"F441",x"EC62",x"F462",x"F482",x"F4A3",x"F4E3",x"F503",x"FCE4",
									 x"FD04",x"FD24",x"FD24",x"FD44",x"FD44",x"FD44",x"FD44",x"FD64",x"FD65",x"FD65",
									 x"FD85",x"FD85",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDC6",
									 x"FDC6",x"FDC6",x"FDC6",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC6",
									 x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",
									 x"FDC6",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDA5",x"FDC5",x"FDA5",
									 x"FDA5",x"FDA5",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",
									 x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",x"FD64",x"FD64",
									 x"FD64",x"FD44",x"FD44",x"FD23",x"FD23",x"F503",x"F503",x"F4E3",x"FCE3",x"FCE3",
									 x"FCC2",x"FCA2",x"FC82",x"FC82",x"F443",x"F443",x"F443",x"F486",x"E4EA",x"E52D",
									 x"E5B2",x"E635",x"D658",x"CE59",x"D69A",x"D6DB",x"DEFC",x"E75D",x"F7BE",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",x"FFBD",x"FF9C",x"FF5B",x"FED8",x"F613",
									 x"ED2E",x"ECCA",x"E467",x"EC64",x"F424",x"FC23",x"F443",x"EC63",x"F483",x"F4A3",
									 x"FCC3",x"FCC4",x"FCE4",x"F504",x"F524",x"FD24",x"FD24",x"FD44",x"FD44",x"FD64",
									 x"FD64",x"FD64",x"FD64",x"FD84",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",
									 x"FDA5",x"FDC5",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",
									 x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FDE6",
									 x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE5",x"FDE5",
									 x"FDE5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC4",x"FDC4",x"FDC4",
									 x"FDC4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",
									 x"FDA4",x"FD84",x"FDA4",x"FD84",x"FD84",x"FD84",x"FD84",x"FD64",x"FD64",x"FD63",
									 x"FD64",x"FD43",x"FD23",x"F523",x"F504",x"F504",x"FCE3",x"FCC3",x"FCA3",x"FCA2",
									 x"F483",x"FC82",x"FC83",x"F463",x"EC86",x"E4A8",x"E4EB",x"E54F",x"DDB2",x"DDF5",
									 x"DE57",x"D6B9",x"D6BA",x"DEDB",x"E71C",x"EF5D",x"F79E",x"FFDF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDE",
									 x"FF7C",x"FF19",x"F675",x"EDD1",x"ED4D",x"ECA8",x"EC44",x"EC03",x"EC23",x"F442",
									 x"FC63",x"FC63",x"F484",x"F4A4",x"FCC4",x"F4E3",x"FD03",x"FD04",x"FD04",x"FD24",
									 x"F544",x"FD44",x"FD44",x"FD64",x"FD84",x"FD84",x"FDA4",x"FDA5",x"FDA5",x"FDA5",
									 x"FDA5",x"FDA5",x"FDC5",x"FDA5",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDE6",x"FDE6",
									 x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",
									 x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDC5",x"FDC4",x"FDC4",x"FDC4",x"FDC4",
									 x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",
									 x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD84",x"FD64",x"FD64",x"FD44",
									 x"FD44",x"FD43",x"FD23",x"FD03",x"FD04",x"FD04",x"FCE4",x"FCE3",x"FCC3",x"F4A3",
									 x"F463",x"EC63",x"EC64",x"EC87",x"E4C9",x"E50C",x"E590",x"D615",x"D637",x"D658",
									 x"DE79",x"DEDB",x"E6FC",x"E75D",x"F79E",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"FFBE",x"FF7C",x"FEF9",x"FE55",x"ED4F",x"EC89",
									 x"EC45",x"F423",x"F421",x"FC42",x"F442",x"FC82",x"FC82",x"FCA3",x"F4E3",x"F4E3",
									 x"FCE3",x"F503",x"F523",x"FD24",x"FD44",x"FD44",x"FD64",x"FD64",x"FD85",x"FD85",
									 x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC6",
									 x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FDE6",x"FE05",x"FDE5",x"FDE5",x"FDE5",
									 x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE4",x"FDE4",x"FDE4",x"FDE4",x"FDE4",x"FDE5",
									 x"FDE5",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",
									 x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD84",x"FD63",x"FD63",x"FD63",x"F543",
									 x"F543",x"F524",x"F503",x"F4E3",x"F4E3",x"F4C3",x"F4A2",x"FC82",x"FC62",x"F463",
									 x"F444",x"EC66",x"E4CA",x"DD4F",x"D5B2",x"D616",x"D658",x"D679",x"D69A",x"DEDB",
									 x"E73C",x"EF9E",x"F7DF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFFF",x"FFDF",x"FFFF",x"FF9D",
									 x"FF1A",x"F697",x"EDF3",x"ED4E",x"EC88",x"F445",x"EC23",x"EC42",x"F462",x"F483",
									 x"F483",x"FCA3",x"FCA3",x"FCC3",x"FCE3",x"F503",x"F524",x"FD24",x"F544",x"F544",
									 x"FD64",x"FD64",x"FD85",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",
									 x"FDA5",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE05",x"FE05",x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDE5",x"FDE5",
									 x"FDE5",x"FDE4",x"FDE4",x"FDE4",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE4",x"FDC4",
									 x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FDA4",
									 x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD84",x"FD64",x"FD64",x"FD43",x"FD23",x"F523",
									 x"F503",x"F4E3",x"F4E3",x"F4C3",x"F4C3",x"F482",x"F463",x"EC64",x"ECA7",x"E4CA",
									 x"DD2C",x"DD90",x"D5F4",x"CE57",x"CE98",x"D699",x"DEDB",x"E73C",x"EF5D",x"F7BF",
									 x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFBC",x"FF7B",x"FED6",x"F5F1",x"ED4D",x"E4C9",x"E466",
									 x"EC44",x"F423",x"F443",x"F482",x"FCA3",x"FCC3",x"FCC4",x"FCC4",x"FCE4",x"FD04",
									 x"FD24",x"FD24",x"FD44",x"FD64",x"FD65",x"FD65",x"FD85",x"FD85",x"FD85",x"FDA5",
									 x"FDA5",x"FDA5",x"FDC5",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDE6",x"FDE6",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE05",x"FE05",
									 x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDE5",x"FDE4",x"FDE4",
									 x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE4",x"FDE5",x"FDE5",x"FDE5",x"FDE4",
									 x"FDE4",x"FDE5",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FDA5",x"FDA4",
									 x"FDA4",x"FD84",x"FD84",x"FD64",x"FD64",x"FD44",x"FD44",x"FD23",x"FD03",x"F503",
									 x"FCE3",x"FCC3",x"FCA3",x"F484",x"EC65",x"EC66",x"EC86",x"E4C9",x"DD2D",x"DDB1",
									 x"D615",x"CE17",x"D659",x"D699",x"DEBA",x"E71C",x"EF7D",x"FFBE",x"FFDF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FFDF",x"FFBF",x"FF7C",x"F6D7",
									 x"F612",x"F56E",x"EC88",x"F424",x"EC23",x"EC22",x"F462",x"F463",x"FC83",x"FCA3",
									 x"FCC3",x"FCE4",x"FCE4",x"FD04",x"FD24",x"FD24",x"FD44",x"FD64",x"FD64",x"FD85",
									 x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDC6",x"FDC6",x"FDE6",
									 x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE26",x"FE26",x"FE26",x"FE26",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE06",x"FE06",x"FE05",x"FE25",x"FE25",x"FE25",x"FE05",x"FE05",
									 x"FE05",x"FE05",x"FE05",x"FE05",x"FE04",x"FE04",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE4",x"FDE4",
									 x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC5",x"FDA5",x"FDA4",x"FDA4",x"FD84",
									 x"FD84",x"FD84",x"FD64",x"FD64",x"FD44",x"FD44",x"F523",x"FD03",x"FCE3",x"FCA3",
									 x"FC83",x"F463",x"F463",x"EC64",x"EC66",x"E4C9",x"DD2E",x"D592",x"D5F6",x"D657",
									 x"D679",x"D6BA",x"DEFB",x"E73C",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDF",x"FFDF",x"FF9E",x"FF3B",x"FE76",x"F5B0",x"F52C",x"EC88",x"F424",x"FC02",
									 x"F422",x"F442",x"F462",x"F4A3",x"F4A2",x"FCE3",x"FD03",x"FD04",x"FD24",x"FD44",
									 x"FD44",x"FD64",x"FD64",x"FD64",x"FD84",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDC5",
									 x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE25",x"FE25",x"FE26",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FDE5",x"FDE5",x"FDE5",x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDE4",x"FDC4",
									 x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD84",
									 x"FD64",x"FD64",x"F544",x"FD43",x"FD23",x"FD03",x"FCC2",x"FCA2",x"F4A2",x"F483",
									 x"F463",x"F464",x"EC87",x"E4EB",x"DD50",x"D5D3",x"D616",x"CE79",x"CE9A",x"D6BB",
									 x"E71C",x"EF7D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FF9C",x"FF19",x"FE54",
									 x"F56E",x"EC88",x"EC45",x"EC24",x"F422",x"FC42",x"F463",x"F483",x"F4A3",x"F4E3",
									 x"F4E3",x"F504",x"FD24",x"FD24",x"FD44",x"F544",x"FD64",x"FD65",x"FD85",x"FD85",
									 x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",
									 x"FDE6",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE26",
									 x"FE26",x"FE26",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE47",
									 x"FE27",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE25",x"FE05",
									 x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FE05",x"FE05",x"FDE4",x"FDE4",x"FDC4",x"FDE5",x"FDE5",x"FDC4",x"FDC4",
									 x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FD84",x"FD84",x"F563",x"F563",
									 x"F543",x"FD23",x"FD23",x"FD03",x"FCE3",x"F4C3",x"F483",x"F463",x"EC63",x"EC65",
									 x"E4CA",x"DD2E",x"DDB2",x"D616",x"CE37",x"CE59",x"DEBA",x"E71C",x"EF5D",x"F7BE",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDF",x"FFBE",x"FF7C",x"EEB6",x"E5D1",x"ED2C",x"EC87",x"EC23",x"F442",x"EC42",
									 x"F462",x"F483",x"F4C4",x"F4C4",x"F504",x"F504",x"F524",x"F524",x"FD44",x"FD64",
									 x"FD64",x"FD85",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC6",
									 x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",x"FE06",x"FE06",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",x"FE05",x"FE05",
									 x"FE05",x"FE25",x"FE25",x"FE25",x"FE05",x"FE25",x"FE05",x"FE25",x"FE25",x"FE25",
									 x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FDE5",x"FE05",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDC4",x"FDC4",x"FDC4",
									 x"FDC4",x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD83",x"FD64",x"FD64",x"F544",x"F524",
									 x"FD23",x"FD03",x"FCC3",x"F4A3",x"F483",x"F464",x"EC85",x"E4A8",x"DD0C",x"D571",
									 x"D5D4",x"CDF7",x"D659",x"D699",x"DEDA",x"E73C",x"F79E",x"F7BF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF9D",x"FEF9",x"F675",x"ED6F",
									 x"E4C9",x"EC66",x"EC24",x"EC22",x"EC42",x"F483",x"F4A3",x"F4C3",x"F4E3",x"F4E3",
									 x"F503",x"F524",x"FD44",x"FD44",x"FD64",x"FD85",x"FD85",x"FD85",x"FD85",x"FDA5",
									 x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDC6",x"FDC6",x"FDE6",x"FE06",x"FDE6",
									 x"FE06",x"FE06",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE27",x"FE27",x"FE27",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE48",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE46",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FE05",x"FE05",x"FDE5",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",
									 x"FDA4",x"FDA4",x"FD84",x"FD64",x"FD44",x"FD44",x"FD24",x"FD23",x"F4E3",x"F4C3",
									 x"F4A3",x"F482",x"F483",x"EC64",x"EC87",x"E4EB",x"D54F",x"CDB3",x"CDF7",x"CE38",
									 x"CE59",x"DEBA",x"EEFC",x"EF5D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFBD",x"FEF8",x"FE13",x"F54E",x"EC89",x"EC25",x"F424",x"FC44",x"FC63",
									 x"F483",x"F4A3",x"FCE3",x"F4E3",x"FD04",x"FD24",x"FD24",x"FD44",x"FD64",x"FD85",
									 x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDC5",x"FDC6",
									 x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",x"FE06",x"FE06",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FDE4",x"FDE4",x"FDE4",x"FDE4",x"FDE4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FD84",
									 x"FD64",x"FD64",x"FD44",x"FD44",x"FD23",x"FD03",x"FCE3",x"F4C3",x"F4A2",x"F482",
									 x"EC64",x"E486",x"DCE9",x"DD2D",x"D593",x"D5F7",x"CE58",x"CE79",x"D69A",x"DEFA",
									 x"EF7C",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFBE",x"FF7C",x"F6D6",x"F5D0",x"F4EB",
									 x"F447",x"F404",x"F402",x"F422",x"F463",x"FCA3",x"F4C3",x"F4E3",x"FD04",x"FD04",
									 x"FD24",x"FD44",x"FD44",x"FD64",x"FD65",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",
									 x"FDA5",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",
									 x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE46",x"FE46",x"FE46",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE05",x"FE05",x"FE05",x"FE04",x"FE04",
									 x"FDE4",x"FDE4",x"FDE4",x"FDC4",x"FDC4",x"FDA4",x"FD84",x"FD84",x"FD84",x"FD64",
									 x"FD44",x"FD24",x"FD23",x"FD03",x"FCE2",x"FCA2",x"F482",x"EC82",x"E484",x"E486",
									 x"DCEC",x"D551",x"CDD4",x"C637",x"CE58",x"CE98",x"DEFA",x"EF5C",x"F7BE",x"FFDE",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",
									 x"FF9D",x"FF1A",x"F695",x"ED8F",x"ECA8",x"EC25",x"F403",x"F422",x"F461",x"F482",
									 x"F4A3",x"F4E3",x"F503",x"F504",x"FD24",x"FD24",x"FD44",x"FD64",x"FD84",x"FD85",
									 x"FD85",x"FDA5",x"FDA5",x"FDC5",x"FDC6",x"FDC5",x"FDC6",x"FDE6",x"FDE6",x"FDE6",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE27",
									 x"FE27",x"FE27",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE27",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE46",x"FE26",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE24",x"FE25",x"FE25",x"FE04",x"FE04",x"FE04",x"FE04",x"FE05",x"FDE5",
									 x"FDE5",x"FDC4",x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD64",x"FD44",x"FD23",
									 x"FD03",x"FCE3",x"FCC3",x"F4A2",x"F482",x"F464",x"EC86",x"DCC9",x"D54E",x"D5D3",
									 x"D617",x"CE18",x"CE79",x"DEFA",x"E73C",x"EF9D",x"FFDE",x"FFDF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFBD",x"FF1A",x"F654",x"F56E",x"F488",
									 x"F424",x"F423",x"F443",x"F463",x"F4A2",x"F4C3",x"F4E4",x"F504",x"FD03",x"FD24",
									 x"FD44",x"FD64",x"FD84",x"FD85",x"FDA5",x"FD85",x"FDA5",x"FDC5",x"FDC6",x"FDC6",
									 x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE26",x"FE26",x"FE26",x"FE27",x"FE27",x"FE27",x"FE27",x"FE48",x"FE48",x"FE48",
									 x"FE48",x"FE48",x"FE48",x"FE48",x"FE48",x"FE68",x"FE68",x"FE68",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE46",x"FE46",x"FE46",x"FE26",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE25",
									 x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",x"FE24",x"FE25",x"FE25",
									 x"FE24",x"FE24",x"FE24",x"FE24",x"FE05",x"FE05",x"FE05",x"FDE5",x"FDC4",x"FDC4",
									 x"FDC4",x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD43",x"FD24",x"FD24",x"F4E4",x"F4C2",
									 x"F4A2",x"F463",x"F464",x"EC85",x"E4E8",x"DD2E",x"DD92",x"CDD6",x"CE38",x"CE79",
									 x"D6BA",x"E73C",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFBD",x"FF3A",x"EE34",x"ED2C",x"EC68",x"F404",x"F422",x"F463",x"EC83",x"F4A3",
									 x"F4C3",x"F4E4",x"F4E4",x"FD04",x"FD24",x"FD44",x"FD64",x"FD65",x"FD85",x"FDA5",
									 x"FDA5",x"FDA5",x"FDA5",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE27",x"FE27",x"FE27",x"FE47",x"FE48",x"FE48",
									 x"FE48",x"FE49",x"FE49",x"FE69",x"FE6A",x"FE6A",x"FE6A",x"FE6A",x"FE6A",x"FE69",
									 x"FE69",x"FE89",x"FE89",x"FE89",x"FE68",x"FE68",x"FE68",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE24",x"FE24",x"FE45",x"FE25",x"FE24",x"FE25",x"FE24",x"FE24",
									 x"FE25",x"FE25",x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDC4",x"FDC4",x"FDA4",x"FDA4",
									 x"FDA4",x"FD84",x"F564",x"FD44",x"F524",x"F503",x"F4E3",x"F4A4",x"F484",x"F464",
									 x"EC85",x"E4A9",x"DD0E",x"D592",x"CDF5",x"CE38",x"CE79",x"D6BA",x"E71C",x"F77E",
									 x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",x"F79B",x"F718",x"FDF2",x"ECCB",x"EC66",
									 x"EC24",x"F442",x"F462",x"F483",x"F4A3",x"F4E4",x"F4E4",x"F504",x"F524",x"FD44",
									 x"FD64",x"FD64",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDC6",x"FDC6",x"FDC6",
									 x"FDE6",x"FDE6",x"FE06",x"FE06",x"FDE5",x"FDE5",x"FE26",x"FE06",x"FE27",x"FE48",
									 x"FE48",x"FE49",x"FE6A",x"FE8B",x"FE6B",x"FE8C",x"FE8B",x"FE8C",x"FE6C",x"FE8C",
									 x"FE8C",x"FE8C",x"FE8C",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",
									 x"FE89",x"FE68",x"FE68",x"FE68",x"FE67",x"FE47",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE44",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE24",x"FE25",x"FE25",x"FE25",x"FE05",
									 x"FE05",x"FE05",x"FDE4",x"FDE4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FD84",x"FD84",
									 x"FD44",x"FD44",x"FD23",x"FD03",x"FCC3",x"FCA2",x"F483",x"EC85",x"E4A8",x"DCEC",
									 x"D570",x"CDD4",x"C5F7",x"C638",x"CEBA",x"E71B",x"EF5D",x"F7BE",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",
									 x"FF7B",x"F6B7",x"F612",x"F50C",x"E425",x"EC24",x"F423",x"F442",x"F483",x"F4A3",
									 x"F4C4",x"FD04",x"FD04",x"FD24",x"FD44",x"FD64",x"FD85",x"FD85",x"FD85",x"FDA5",
									 x"FDC5",x"FDC6",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FE06",x"FE27",x"FE48",x"FE69",x"FE6A",x"FE8B",x"FE8B",x"FEAC",x"FEAC",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAD",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FE8B",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE6A",x"FE89",x"FE89",x"FE69",
									 x"FE68",x"FE68",x"FE68",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",
									 x"FE46",x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE25",x"FE45",x"FE45",x"FE25",x"FE25",x"FE25",x"FE05",x"FE05",x"FE04",
									 x"FDE4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD64",x"FD44",x"FD23",
									 x"FD03",x"FCC2",x"FCA2",x"F483",x"EC65",x"E487",x"DCEB",x"D571",x"CDB4",x"C5F7",
									 x"C658",x"D69A",x"DEFB",x"EF5C",x"FFDE",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFE",x"FFFF",x"FFFF",x"FFFF",x"FF9D",x"FEB7",x"F590",x"F4EB",x"F466",
									 x"EC03",x"F443",x"FC63",x"FC83",x"F4A3",x"F4C4",x"F4E4",x"FD04",x"FD24",x"FD24",
									 x"FD44",x"FD85",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDC5",x"FDC6",x"FDC6",x"FDC5",
									 x"FDE5",x"FDE6",x"FE06",x"FE26",x"FE26",x"FE27",x"FE28",x"FE49",x"FE6A",x"FE8C",
									 x"FEAD",x"FEAD",x"FEAD",x"FEAD",x"FECE",x"FEAD",x"FEAD",x"FEAD",x"FEAD",x"FEAD",
									 x"FECD",x"FECD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8C",x"FE8B",
									 x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE6A",x"FE69",x"FE69",x"FE69",x"FE68",x"FE67",
									 x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",
									 x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE26",x"FE26",x"FE26",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE65",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE25",x"FE25",x"FE25",x"FE24",x"FE25",x"FE05",x"FE04",x"FDE4",x"FDE4",x"FDC4",
									 x"FDC4",x"FDA4",x"FDA4",x"FD84",x"FD64",x"FD44",x"FD23",x"FD03",x"FCC2",x"FCA2",
									 x"FCA3",x"F484",x"EC86",x"ECEB",x"DD51",x"CDB4",x"C616",x"CE38",x"D679",x"DEDB",
									 x"EF7D",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",x"FFBD",
									 x"FF5C",x"FED7",x"FD8F",x"EC68",x"EC25",x"F422",x"F421",x"F462",x"FCA3",x"FCC3",
									 x"FCE4",x"F504",x"F504",x"FD24",x"FD45",x"FD44",x"FD64",x"FD85",x"FDA5",x"FDA5",
									 x"FDA5",x"FDC6",x"FDC6",x"FDE6",x"FDC6",x"FDE6",x"FE06",x"FE07",x"FE28",x"FE48",
									 x"FE49",x"FE6B",x"FE8C",x"FE8D",x"FEAF",x"FECF",x"FEB0",x"FECF",x"FECF",x"FECF",
									 x"FECE",x"FECE",x"FEAE",x"FEAD",x"FEAD",x"FEAD",x"FECD",x"FEAD",x"FEAC",x"FEAC",
									 x"FEAB",x"FE8B",x"FE8B",x"FE8C",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE6B",x"FE6A",
									 x"FE8A",x"FE6A",x"FE6A",x"FE69",x"FE68",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE46",x"FE46",x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE44",
									 x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE24",
									 x"FE25",x"FE25",x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDE4",x"FDC4",x"FDC4",x"FDA4",
									 x"FD84",x"FD84",x"F564",x"F544",x"F504",x"F4E3",x"F4C3",x"F4A3",x"F464",x"F487",
									 x"E4CB",x"D52F",x"CDB3",x"CDD6",x"CE18",x"D679",x"DEFC",x"E75D",x"EF9E",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FF5A",x"F696",x"F5B0",x"ECA8",x"EC04",
									 x"EC23",x"F442",x"F462",x"F4A2",x"F4C3",x"FD04",x"FD24",x"F524",x"FD24",x"FD44",
									 x"FD65",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDC5",x"FDC6",x"FDE6",x"FDE6",x"FDE6",
									 x"FDE6",x"FE07",x"FE28",x"FE29",x"FE4A",x"FE6C",x"FE8D",x"FEAF",x"FEAF",x"FED0",
									 x"FED1",x"FED0",x"FEB0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FEAE",x"FEAE",
									 x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FE8B",
									 x"FEAB",x"FE8B",x"FEAB",x"FE8B",x"FE6A",x"FE6A",x"FE6A",x"FE6A",x"FE69",x"FE69",
									 x"FE68",x"FE68",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE26",
									 x"FE26",x"FE26",x"FE25",x"FE25",x"FE45",x"FE25",x"FE25",x"FE25",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE44",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",
									 x"FE05",x"FE05",x"FE04",x"FDE4",x"FDE4",x"FDC4",x"FDA4",x"FDA4",x"F584",x"F564",
									 x"F544",x"F524",x"F4E3",x"F4C3",x"F4A3",x"F464",x"EC66",x"E4A9",x"DD4E",x"D5B3",
									 x"CDF6",x"CE17",x"D69A",x"DF1C",x"E75D",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",
									 x"FF7C",x"FEB6",x"ED8F",x"F4CA",x"EC45",x"EC22",x"EC42",x"EC63",x"F4A3",x"F4E3",
									 x"F4E3",x"F504",x"F524",x"F524",x"FD44",x"FD64",x"FD85",x"FD85",x"FDA5",x"FDC5",
									 x"FDA5",x"FDC5",x"FDC6",x"FDE6",x"FDE6",x"FE06",x"FE27",x"FE28",x"FE4A",x"FE6C",
									 x"FE8E",x"FEAF",x"FED0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FEAF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FEAE",x"FEAE",x"FEAE",x"FEAD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAB",x"FEAB",x"FEAB",x"FE8B",x"FE8B",
									 x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE69",x"FE68",x"FE68",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE25",
									 x"FE44",x"FE44",x"FE45",x"FE65",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE25",x"FE25",x"FE25",x"FE05",x"FE04",
									 x"FDE4",x"FDC4",x"FDC4",x"FDA4",x"FD84",x"FD84",x"FD64",x"FD44",x"FD03",x"F4E3",
									 x"F4C3",x"F483",x"F464",x"EC65",x"DCCA",x"D550",x"CDB4",x"CDF6",x"CE39",x"CE9A",
									 x"DEFC",x"EF7D",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FF7D",x"FEB7",x"F56E",x"EC88",x"EC45",
									 x"EC23",x"F443",x"F463",x"F4A4",x"F4C4",x"F4E4",x"FD04",x"FD24",x"FD44",x"FD44",
									 x"FD64",x"FD64",x"FD85",x"FDA5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC6",x"FDE7",
									 x"FE08",x"FE29",x"FE4A",x"FE6C",x"FE8E",x"FEAF",x"FED0",x"FED0",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",
									 x"FEAE",x"FEAD",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE8A",
									 x"FE8A",x"FE89",x"FE69",x"FE69",x"FE68",x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",
									 x"FE46",x"FE26",x"FE26",x"FE26",x"FE45",x"FE45",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE24",x"FE24",x"FE24",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE44",x"FE44",x"FE45",x"FE65",x"FE65",x"FE85",
									 x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE45",
									 x"FE45",x"FE45",x"FE25",x"FE25",x"FE04",x"FE04",x"FE04",x"FDE4",x"FDC4",x"FDC4",
									 x"FDA4",x"FDA4",x"FD84",x"FD64",x"FD44",x"F523",x"F503",x"F4C2",x"F483",x"F464",
									 x"E487",x"DCEB",x"DD4E",x"D593",x"CDF7",x"C638",x"CE7A",x"E6FC",x"EF7D",x"F7BE",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",
									 x"FF1A",x"FE76",x"F590",x"E447",x"EC24",x"EC23",x"F443",x"FC83",x"F4A2",x"F4C3",
									 x"FCE4",x"FD04",x"FD24",x"FD44",x"FD44",x"FD65",x"FD85",x"FD86",x"FDA6",x"FDC6",
									 x"FDC6",x"FDC6",x"FDC5",x"FDC5",x"FDE7",x"FE29",x"FE4B",x"FE6D",x"FEAE",x"FED0",
									 x"FED1",x"FED2",x"FED2",x"FED1",x"FEF1",x"FED0",x"FED0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FEAE",x"FECE",x"FEAD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",
									 x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE69",x"FE69",
									 x"FE68",x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE26",x"FE26",x"FE25",
									 x"FE45",x"FE46",x"FE46",x"FE46",x"FE45",x"FE45",x"FE45",x"FE45",x"FE66",x"FE66",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",
									 x"FE65",x"FE85",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",
									 x"FE25",x"FE25",x"FE05",x"FE05",x"FDE5",x"FE05",x"FDE5",x"FDC4",x"FDA4",x"FDA4",
									 x"FD64",x"FD44",x"F543",x"F502",x"F4C2",x"F4A3",x"EC84",x"E486",x"E4A9",x"DD0D",
									 x"CD93",x"C5D6",x"C5F7",x"D659",x"DEDB",x"E75C",x"F7BE",x"FFDF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FF7B",x"F613",x"ED2D",x"EC88",x"EBE4",
									 x"F423",x"F442",x"FC82",x"FCA2",x"F4C3",x"F4E3",x"FD04",x"FD24",x"FD45",x"FD65",
									 x"FD85",x"FD85",x"FDA5",x"FDA6",x"FDA6",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FE07",
									 x"FE4A",x"FE8C",x"FEAF",x"FED1",x"FED2",x"FEF3",x"FEF3",x"FED3",x"FED2",x"FED1",
									 x"FED0",x"FED0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FEEF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",
									 x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE69",x"FE69",x"FE68",x"FE48",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE46",x"FE46",x"FE26",x"FE25",x"FE45",x"FE46",x"FE46",x"FE46",x"FE65",
									 x"FE84",x"FE84",x"FEA5",x"FEA6",x"FEC6",x"FEC6",x"FEC6",x"FEA5",x"FE85",x"FE85",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE44",x"FE45",x"FE45",x"FE45",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",
									 x"FE05",x"FE05",x"FDE5",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD64",x"F563",x"F543",
									 x"FD02",x"FCC2",x"FCA3",x"F484",x"F464",x"E488",x"D52E",x"CDB3",x"C5D6",x"C617",
									 x"CE79",x"DEDA",x"EF5D",x"F7BF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",
									 x"FFBD",x"FEF8",x"F58F",x"F4A8",x"EC45",x"EC03",x"F422",x"F462",x"F483",x"F4C3",
									 x"F4E4",x"FD04",x"FD25",x"FD44",x"FD65",x"FD85",x"FD85",x"FDA5",x"FDC5",x"FDC5",
									 x"FDC5",x"FDC5",x"FDE6",x"FE07",x"FE28",x"F64A",x"FE8D",x"FED0",x"FED2",x"FEF3",
									 x"FEF3",x"FEF3",x"FEF2",x"FEF2",x"FED1",x"FED0",x"FED0",x"FED0",x"FED0",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",
									 x"FE69",x"FE69",x"FE68",x"FE68",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE46",
									 x"FE45",x"FE45",x"FE46",x"FE46",x"FE65",x"FE64",x"FE85",x"FE65",x"FE85",x"FE86",
									 x"FEA6",x"FEC6",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FEA5",x"FE84",
									 x"FE84",x"FE84",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",x"FE05",x"FE04",x"FDE4",
									 x"FDE4",x"FDC4",x"FDA4",x"FD84",x"F584",x"F544",x"F523",x"FCE3",x"FCA3",x"FC63",
									 x"FC43",x"EC65",x"DCEB",x"D590",x"CDB3",x"C5D6",x"C638",x"CE99",x"E71B",x"EF7E",
									 x"F7BF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FF7C",x"FEF8",x"EDD1",x"ECA9",x"EC24",
									 x"EC23",x"F463",x"F483",x"F4A3",x"F4C4",x"F504",x"F504",x"FD25",x"FD45",x"FD64",
									 x"FD85",x"FD85",x"FDA5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDE6",x"F608",x"FE4B",
									 x"FE8D",x"FEAF",x"FED1",x"FEF2",x"FEF3",x"FEF3",x"FEF2",x"FEF2",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",
									 x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE69",x"FE68",x"FE68",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE46",x"FE26",x"FE46",x"FE25",x"FE45",x"FE46",x"FE26",
									 x"F605",x"E5A5",x"D505",x"CCE5",x"CCE5",x"CD05",x"D565",x"DD85",x"E5C5",x"E605",
									 x"EE45",x"F666",x"FEA6",x"FEC6",x"FEC6",x"FEE6",x"FEE5",x"FEC5",x"FEA5",x"FE85",
									 x"FEA5",x"F664",x"F664",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE84",x"FE84",x"FE84",x"FE85",x"FE85",x"FE85",x"FE65",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE65",
									 x"FE45",x"FE45",x"FE45",x"FE25",x"FE05",x"FE04",x"FDE4",x"FDE4",x"FDC4",x"FDA4",
									 x"FD84",x"F564",x"F564",x"F523",x"FCE3",x"FCA3",x"FC83",x"F484",x"E4A7",x"DCEB",
									 x"D52E",x"CD93",x"C5F6",x"C638",x"D69A",x"E71C",x"EF7E",x"F7BE",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",
									 x"FF7C",x"F6B7",x"F5D1",x"ECA9",x"EC04",x"F402",x"F422",x"FCA3",x"F4C3",x"F4E3",
									 x"F504",x"F524",x"F524",x"FD44",x"FD64",x"FD65",x"FD85",x"FDA5",x"FDA5",x"FDC5",
									 x"FDE5",x"FDC5",x"FDE6",x"FE29",x"FE6C",x"FED0",x"FEF2",x"FEF2",x"FEF3",x"FF14",
									 x"FEF3",x"FEF2",x"FEF1",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECE",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",
									 x"FE8A",x"FE89",x"FE89",x"FE89",x"FE68",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE47",x"FE46",x"FE24",x"FE45",x"FE26",x"E584",x"C483",x"A362",x"8261",x"7A42",
									 x"7A41",x"8261",x"8AC1",x"9321",x"9B82",x"AC02",x"B443",x"BCA3",x"CD24",x"D584",
									 x"DDC4",x"E624",x"EE64",x"EEA4",x"F6A5",x"FEE5",x"FF06",x"FEE5",x"FEC5",x"FEA5",
									 x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE84",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",
									 x"FE25",x"FE04",x"FE04",x"FDE4",x"FDE4",x"FDC4",x"FDA4",x"FD83",x"FD83",x"F564",
									 x"F524",x"F4E3",x"FCC3",x"F4A3",x"EC84",x"EC66",x"E4AA",x"DD50",x"CDB4",x"BDF7",
									 x"C618",x"D69A",x"E71C",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFFF",x"FFBE",x"FEF9",x"F5F2",x"F4EB",x"EC25",
									 x"F402",x"FC42",x"F442",x"FCC3",x"F4C3",x"F4E3",x"F504",x"FD24",x"FD44",x"FD64",
									 x"FD84",x"F585",x"FD85",x"FD85",x"FDA4",x"FDC5",x"FDC5",x"FDE6",x"FE29",x"FE6D",
									 x"FED0",x"FF12",x"FF13",x"FF14",x"FF13",x"FEF3",x"FEF2",x"FEF2",x"FEF1",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",
									 x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE69",
									 x"FE68",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE47",x"FE46",x"FE24",x"FE65",
									 x"F606",x"CCA5",x"9302",x"6180",x"50E0",x"48A0",x"4880",x"48A0",x"58E0",x"6140",
									 x"69A0",x"7A41",x"8AA1",x"9302",x"A382",x"AC03",x"B463",x"C4E3",x"D584",x"DDE5",
									 x"EE65",x"F6E6",x"FF46",x"FF46",x"FF26",x"FF06",x"FEC6",x"FEA5",x"F685",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FEA4",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE24",x"FE04",
									 x"FDE4",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD64",x"FD44",x"F503",x"FD03",x"FCC3",
									 x"F4A3",x"F464",x"EC46",x"E4EC",x"D572",x"C5D5",x"BDF6",x"C659",x"D6BB",x"DF1C",
									 x"EFBE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDE",x"FF5A",x"F633",x"ED0C",x"EC67",x"EC04",x"F422",x"FC63",x"F463",x"F4C3",
									 x"F4E3",x"F504",x"FD24",x"FD44",x"FD64",x"FD64",x"FD85",x"FDA5",x"FDA5",x"FDA4",
									 x"FDA5",x"FDC7",x"FDE8",x"FE2B",x"FE6D",x"FED1",x"FEF3",x"FF14",x"FF14",x"FEF4",
									 x"FEF3",x"FEF3",x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8B",x"FE8A",
									 x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE69",x"FE68",x"FE68",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE47",x"FE47",x"FE45",x"FE44",x"E565",x"A382",x"69E1",x"48A0",
									 x"4060",x"4880",x"4880",x"50A0",x"58E0",x"6100",x"6140",x"6960",x"71A0",x"71E0",
									 x"79E1",x"7A21",x"7A40",x"82A1",x"9B62",x"A3E3",x"B483",x"C544",x"D605",x"DE64",
									 x"EEC4",x"F725",x"FF45",x"FF46",x"FF05",x"FEC5",x"FEA5",x"FE85",x"FE64",x"FE65",
									 x"FE65",x"FE66",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE04",x"FE04",x"FDE4",x"FDC4",x"FDC4",
									 x"FDA4",x"FD84",x"FD64",x"FD23",x"FD23",x"FD03",x"F4C2",x"FC82",x"F464",x"E4A9",
									 x"DD0D",x"D592",x"C5D5",x"C617",x"CE39",x"D6BA",x"E75C",x"F7BE",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FF3A",x"FE54",x"ED0B",x"EC46",
									 x"EC04",x"F443",x"FC62",x"FCA3",x"F4C3",x"F4E4",x"F524",x"FD24",x"FD45",x"FD65",
									 x"FD64",x"FD84",x"FDA5",x"FDA5",x"FDC4",x"FDC4",x"FDE7",x"FE0A",x"FE6D",x"FED0",
									 x"FEF2",x"FF14",x"FF15",x"FF15",x"FF14",x"FF13",x"FEF3",x"FEF3",x"FEF2",x"FEF2",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE8A",
									 x"FE89",x"FE69",x"FE68",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE47",
									 x"FE46",x"FE25",x"CCC4",x"8280",x"5100",x"3840",x"4881",x"58E1",x"6101",x"6921",
									 x"6941",x"6940",x"6940",x"6920",x"6920",x"6120",x"6100",x"60E0",x"58E0",x"5900",
									 x"6960",x"71E1",x"7A40",x"82C2",x"9382",x"9C01",x"ACE1",x"CDC3",x"E664",x"EEC5",
									 x"F705",x"FF05",x"FF05",x"FF04",x"FEE4",x"FEC5",x"FEA5",x"FE85",x"FE66",x"FE66",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",x"FE45",
									 x"FE45",x"FE25",x"FE25",x"FE05",x"FDE5",x"FDC5",x"FDC4",x"FDA4",x"FD84",x"FD64",
									 x"F543",x"F522",x"F502",x"FCC2",x"FCA3",x"EC85",x"E488",x"DD0D",x"D5B2",x"C5F6",
									 x"C5F8",x"CE39",x"DEDA",x"EF5C",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FF5C",x"FE96",x"FD6E",x"EC26",x"F3E3",x"F423",x"F462",x"F482",x"FCC3",
									 x"F4E4",x"F504",x"F524",x"F524",x"FD45",x"FD65",x"FD85",x"FDA5",x"FDA5",x"FDC4",
									 x"FDC4",x"FE06",x"FE49",x"FE8D",x"FED1",x"FF13",x"FF34",x"FF34",x"FF34",x"FF13",
									 x"FF14",x"FF13",x"FF13",x"FEF3",x"FEF2",x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",
									 x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE69",x"FE68",x"FE67",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE46",x"FE46",x"FE26",x"C4A4",x"7A60",
									 x"5100",x"4060",x"50C1",x"6120",x"6120",x"7140",x"7140",x"7161",x"7981",x"7161",
									 x"7961",x"7161",x"7180",x"7181",x"7181",x"6961",x"6961",x"6961",x"6940",x"6960",
									 x"6180",x"61E0",x"7AA0",x"9BA2",x"AC62",x"BD04",x"D5E5",x"EEC6",x"FF46",x"FF85",
									 x"FF65",x"FF25",x"FEE4",x"FEA4",x"FE84",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",x"FE45",x"FE25",
									 x"FE05",x"FDE5",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"F583",x"F543",x"FD03",x"FCE3",
									 x"F4C2",x"F463",x"F466",x"E4A9",x"D56F",x"CDB5",x"C5D7",x"BDF8",x"CE9A",x"DEFB",
									 x"EF5D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FED8",x"FDB1",x"FCA9",
									 x"EBE3",x"F402",x"F443",x"F483",x"F4C2",x"FCE3",x"F4E4",x"FD24",x"FD44",x"FD45",
									 x"FD65",x"FD85",x"F584",x"FDA4",x"FDC5",x"FDC5",x"FE07",x"FE49",x"FE8D",x"FEF1",
									 x"FF13",x"FF35",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FEF3",x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",
									 x"FE8A",x"FE89",x"FE69",x"FE69",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",
									 x"FE46",x"FE46",x"FE66",x"FE46",x"C4C4",x"8280",x"5100",x"4080",x"50C0",x"6120",
									 x"6940",x"7160",x"7160",x"7981",x"79A1",x"79A1",x"7981",x"81C1",x"79C0",x"79C0",
									 x"79C0",x"71C1",x"6980",x"6960",x"6960",x"6140",x"5920",x"5940",x"69C1",x"7A42",
									 x"82C3",x"8B43",x"AC65",x"CD65",x"DE46",x"EEC6",x"FF26",x"FF66",x"FF45",x"FF05",
									 x"FEC4",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FEA5",x"FE85",x"FE85",
									 x"FE85",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",x"FE25",x"FE25",x"FE05",x"FE04",x"FDE4",
									 x"FDC4",x"FDA4",x"FDA4",x"FD64",x"FD24",x"F503",x"F502",x"F4A3",x"FC64",x"EC86",
									 x"DCEA",x"D570",x"CDB5",x"C5D7",x"C638",x"D6BA",x"E71C",x"EF7D",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFDE",x"F739",x"EDF2",x"ECCA",x"F424",x"F402",x"F462",x"F483",x"F4C3",
									 x"F4E3",x"FD04",x"FD05",x"FD24",x"FD44",x"FD65",x"FD85",x"FDA5",x"FDA5",x"FDA5",
									 x"FDC5",x"FDE7",x"FE2B",x"FE8F",x"FEF2",x"FF34",x"FF35",x"FF15",x"FF35",x"FF34",
									 x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FEF3",x"FEF2",x"FEF2",x"FEF2",
									 x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",
									 x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE69",x"FE69",
									 x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE46",x"FE46",x"FE46",x"FE26",x"FE26",x"FE46",x"FE46",x"FE46",x"FE65",x"FE45",
									 x"CD04",x"8AE1",x"6141",x"4060",x"50C0",x"6141",x"6960",x"7161",x"7160",x"79A1",
									 x"79A0",x"81C1",x"79A0",x"81E0",x"79C0",x"79C0",x"71C0",x"71C1",x"71A1",x"69A1",
									 x"69A0",x"61A0",x"61A0",x"61A0",x"6180",x"6160",x"5940",x"6180",x"7240",x"8B01",
									 x"9BE2",x"B4A4",x"D5E4",x"EEA6",x"F727",x"FF47",x"FF26",x"FEE5",x"FEA5",x"FEA5",
									 x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",
									 x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",
									 x"FE65",x"FE45",x"FE25",x"FE25",x"FE04",x"FE04",x"FDE4",x"FDC4",x"FDC4",x"FD84",
									 x"FD44",x"F543",x"F543",x"F4E2",x"FC62",x"FC63",x"E486",x"DCEB",x"D571",x"CDB4",
									 x"C5F6",x"CE59",x"D6BA",x"E73C",x"F79E",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",x"FFFF",x"F7DE",x"FF5B",x"F633",x"E50B",
									 x"EC45",x"F3E2",x"FC22",x"FC83",x"F4A3",x"FCE4",x"FD04",x"FD24",x"FD24",x"FD65",
									 x"FD65",x"FD84",x"FDA4",x"FDC5",x"FDA5",x"FDC5",x"FDE8",x"FE4C",x"FEB0",x"FEF3",
									 x"FF35",x"FF36",x"FF16",x"FF15",x"FF15",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FEF2",x"FEF2",x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",
									 x"FE8A",x"FE8A",x"FE89",x"FE6A",x"FE69",x"FE48",x"FE68",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE26",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE45",x"FE66",x"E585",x"A382",x"6981",x"4060",
									 x"50C1",x"6141",x"6940",x"7160",x"7980",x"79A0",x"79C0",x"81C0",x"81A0",x"79A0",
									 x"71A0",x"7180",x"7161",x"6960",x"6160",x"6160",x"61A0",x"61A0",x"61C0",x"61A0",
									 x"6180",x"6180",x"6180",x"6160",x"6180",x"69C1",x"7200",x"8261",x"9BA1",x"B4A3",
									 x"C563",x"E685",x"F746",x"FF67",x"FF46",x"FF06",x"FEE6",x"FEC6",x"FEA5",x"FEA5",
									 x"FEA5",x"FEA5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",
									 x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",
									 x"FE24",x"FE05",x"FE04",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD63",x"F543",x"F503",
									 x"FCC2",x"FC82",x"EC84",x"E4A7",x"DD0C",x"CD92",x"C5D5",x"BDF7",x"C658",x"D6DA",
									 x"EF3C",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFDF",x"FF7C",x"FEB6",x"F54E",x"E468",x"EC23",x"F422",x"FC43",x"FC83",
									 x"F4A3",x"FCE4",x"FD04",x"FD24",x"FD44",x"FD65",x"FD85",x"FD85",x"FD84",x"FDA4",
									 x"F5A5",x"FDE7",x"FE4B",x"FEB0",x"FF13",x"FF35",x"FF56",x"FF16",x"FF15",x"FF15",
									 x"FF15",x"FF14",x"FF34",x"FF33",x"FF33",x"FF13",x"FF13",x"FF13",x"FEF2",x"FEF2",
									 x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE6A",
									 x"FE69",x"FE48",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE46",x"FE26",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE45",x"FE66",x"EDC6",x"B402",x"71E1",x"4060",x"50A0",x"6141",x"6960",x"7160",
									 x"7980",x"79A0",x"81C0",x"81A0",x"79A1",x"71A1",x"71C2",x"71C3",x"69C3",x"69C3",
									 x"6181",x"59A1",x"5980",x"5180",x"5980",x"5960",x"5980",x"6181",x"61C0",x"61A0",
									 x"61A1",x"6180",x"6180",x"69A0",x"7A40",x"8B21",x"A3E2",x"C544",x"E686",x"EF06",
									 x"F746",x"F725",x"F705",x"FF05",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",
									 x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",
									 x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE05",x"FE04",
									 x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD44",x"F524",x"FCE3",x"FCC2",x"F4A3",x"EC85",
									 x"E4A8",x"D52E",x"CDB4",x"C5D7",x"BDF7",x"CE79",x"E6FB",x"EF5D",x"F7BE",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FEB7",x"FDB0",
									 x"F4A9",x"EC04",x"F442",x"F442",x"F483",x"FCC4",x"FCC3",x"FD04",x"FD24",x"FD44",
									 x"FD45",x"FD85",x"FD85",x"FD85",x"FD84",x"FDA4",x"F5E7",x"F64C",x"FED0",x"FF13",
									 x"FF35",x"FF56",x"FF36",x"FF15",x"FF15",x"FF15",x"FF14",x"FF34",x"FF34",x"FF33",
									 x"FF33",x"FF13",x"FF13",x"FF13",x"FEF2",x"FEF2",x"FEF2",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",
									 x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE89",x"FE69",x"FE68",x"FE68",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",
									 x"FE26",x"FE46",x"FE46",x"FE46",x"FE26",x"FE46",x"FE45",x"FE86",x"F605",x"C4A3",
									 x"8281",x"50E0",x"50C0",x"6101",x"6940",x"7160",x"7981",x"79A0",x"79C0",x"7980",
									 x"81E2",x"8265",x"8B09",x"936B",x"938C",x"8B6B",x"7AE8",x"6A65",x"59E3",x"4981",
									 x"4940",x"4920",x"5140",x"5981",x"61C0",x"61E0",x"69C1",x"69E1",x"69C0",x"69C0",
									 x"71C0",x"7A01",x"7A20",x"9342",x"AC62",x"C543",x"DE85",x"F767",x"FFA7",x"FF65",
									 x"FF05",x"F6E5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",
									 x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE65",x"FE65",x"FE45",x"FE25",x"FE04",x"FDE4",x"FDE4",x"FDA4",x"FDA4",
									 x"FD84",x"FD44",x"FD24",x"F503",x"F4C3",x"F482",x"F465",x"DCCA",x"D550",x"CDD6",
									 x"BDF7",x"C638",x"D69B",x"E6FB",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFDF",x"FF3A",x"F5B1",x"F4AA",x"FC25",x"F403",x"F462",x"F482",
									 x"F4C3",x"FCC4",x"FCE4",x"FD04",x"FD25",x"FD45",x"FD65",x"FD85",x"FD85",x"FD85",
									 x"FDA5",x"FDE7",x"FE2B",x"FEB0",x"FF34",x"FF56",x"FF56",x"FF56",x"FF35",x"FF35",
									 x"FF14",x"FF14",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",
									 x"FE89",x"FE89",x"FE68",x"FE68",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE26",x"FE46",x"FE46",x"FE46",
									 x"FE26",x"FE46",x"FE46",x"FE85",x"FE46",x"D524",x"9B42",x"6980",x"58E1",x"5901",
									 x"6940",x"7181",x"7981",x"79A0",x"79A0",x"79A0",x"8265",x"936A",x"A491",x"B533",
									 x"B554",x"AD33",x"9CB0",x"8C0D",x"838A",x"6AC7",x"5A24",x"51E3",x"4961",x"4960",
									 x"5180",x"59C0",x"61E0",x"69E1",x"6A01",x"7201",x"69C0",x"71C0",x"71A1",x"7A01",
									 x"8280",x"9341",x"AC83",x"D606",x"E6A6",x"FF45",x"FF65",x"FF45",x"FF05",x"FEE5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEC5",x"FEC5",x"FEC5",
									 x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",
									 x"FE45",x"FE25",x"FE04",x"FDE4",x"FDC4",x"FDC4",x"FDA4",x"FD64",x"F544",x"F523",
									 x"F4E2",x"FCA2",x"FC63",x"EC86",x"DCEC",x"D593",x"C5D5",x"BDF7",x"CE59",x"D69A",
									 x"E71B",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FFDE",x"FF9C",x"FE95",
									 x"F4EB",x"F446",x"F403",x"F443",x"FC82",x"F4A3",x"FCE4",x"F504",x"FD04",x"FD04",
									 x"FD25",x"FD65",x"FD65",x"FD85",x"FD85",x"FD86",x"FDC7",x"FE4B",x"FE8F",x"FF14",
									 x"FF56",x"FF36",x"FF56",x"FF36",x"FF35",x"FF35",x"FF14",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FEF2",x"FEF2",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",
									 x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE68",x"FE67",
									 x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE45",x"FE85",
									 x"FE65",x"E584",x"ABE2",x"7A21",x"5900",x"58E0",x"6941",x"7181",x"7980",x"7180",
									 x"79A0",x"79C2",x"8AE7",x"A44E",x"B595",x"BE18",x"BE38",x"BE17",x"B5B5",x"B553",
									 x"AD12",x"9CB0",x"8BEC",x"7B6A",x"5A45",x"4181",x"4960",x"4980",x"59A0",x"61E0",
									 x"6A01",x"7201",x"7200",x"7A01",x"7A01",x"81E1",x"7A01",x"7A40",x"8B01",x"A403",
									 x"BD04",x"E645",x"FF47",x"FF86",x"FF66",x"F705",x"F6E5",x"FEE5",x"FEC5",x"FEA5",
									 x"FEA5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",
									 x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE25",x"FE25",x"FE04",
									 x"FDE4",x"FDC4",x"FDA4",x"FD83",x"FD63",x"F543",x"F503",x"FCC2",x"FC82",x"EC64",
									 x"E4C8",x"E52E",x"CD92",x"C5F6",x"C5F8",x"CE59",x"DEDA",x"EF7D",x"F7BE",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFDE",x"FFBD",x"FF3A",x"F5AF",x"EC66",x"EC04",x"EC43",x"F483",
									 x"FCA3",x"FCC3",x"FCE4",x"FD04",x"FD24",x"FD25",x"FD45",x"FD65",x"FD85",x"FD85",
									 x"FD85",x"FDA6",x"FE0A",x"FECF",x"FF13",x"FF36",x"FF36",x"FF36",x"FF35",x"FF35",
									 x"FF35",x"FF15",x"FF15",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF1",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",
									 x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE68",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE26",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE45",x"FE26",x"FE45",x"FE65",x"FE66",x"EDE5",x"C463",x"8AA2",
									 x"50E0",x"50C0",x"6120",x"7181",x"7980",x"7180",x"79A0",x"7A02",x"8B29",x"A490",
									 x"B5D7",x"BE18",x"B618",x"BE18",x"BDF7",x"BDD6",x"BDD6",x"BDB6",x"AD33",x"A4B0",
									 x"83AB",x"5A45",x"4961",x"4160",x"51A0",x"59C0",x"61C0",x"61C0",x"7221",x"7A21",
									 x"8221",x"8221",x"8220",x"8220",x"8260",x"8AC1",x"9B82",x"BCC4",x"DE26",x"EEC6",
									 x"F746",x"FF66",x"FF46",x"FF26",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE65",x"FE65",x"FE45",x"FE25",x"FE05",x"FDE4",x"FDE4",x"FDC4",x"FDA3",
									 x"FD83",x"FD43",x"F524",x"F4E3",x"F4C3",x"F483",x"EC85",x"E4CA",x"D54F",x"CDD5",
									 x"C5D7",x"C618",x"D679",x"E71C",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"FEF9",
									 x"FE33",x"ECCA",x"EC24",x"F422",x"F442",x"F483",x"F4A3",x"FCE4",x"FD04",x"FD24",
									 x"FD44",x"FD45",x"FD46",x"FD85",x"FDA4",x"F5C5",x"FDC7",x"FE0A",x"FE90",x"FF15",
									 x"FF36",x"FF36",x"FF36",x"FF36",x"FF36",x"FF35",x"FF35",x"FF15",x"FF14",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FF11",x"FEF0",x"FEF0",x"FED0",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FE8C",x"FEAB",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE69",
									 x"FE68",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE26",x"FE26",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE25",
									 x"FE25",x"FE65",x"FE85",x"F645",x"D523",x"A364",x"6100",x"50A0",x"6120",x"6980",
									 x"7180",x"7160",x"71A0",x"79E3",x"932A",x"ACB1",x"BDD7",x"BDF9",x"B5F8",x"BDF7",
									 x"BE17",x"C618",x"C639",x"C639",x"CE38",x"CE37",x"BD95",x"8C0E",x"5A86",x"51E3",
									 x"4940",x"5180",x"61C0",x"61E1",x"7241",x"7A41",x"8261",x"8A61",x"8A61",x"8A41",
									 x"8240",x"8220",x"8240",x"92E0",x"B443",x"CD44",x"DE65",x"F746",x"FF86",x"FF85",
									 x"FF45",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEC5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",
									 x"FE25",x"FE25",x"FE05",x"FDE4",x"FDE4",x"FDC4",x"FDA4",x"FD64",x"F544",x"F523",
									 x"F4E3",x"F4A3",x"F484",x"EC67",x"DCEA",x"CD91",x"C5B7",x"BDD9",x"C638",x"D6DB",
									 x"E73D",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"F7DF",x"FFFF",x"FFDE",x"FF5B",x"EE34",x"F54D",x"EC26",x"EC03",x"F422",
									 x"F462",x"F4A4",x"F4C4",x"FD04",x"FD24",x"FD44",x"FD64",x"FD65",x"FD65",x"FD84",
									 x"FDA4",x"F5E6",x"FE2A",x"FE8E",x"FEF3",x"FF37",x"FF57",x"FF36",x"FF35",x"FF36",
									 x"FF36",x"FF35",x"FF35",x"FF15",x"FF14",x"FF34",x"FF34",x"FF34",x"FF34",x"FF33",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FF11",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAB",x"FE8B",x"FE8B",
									 x"FE8B",x"FE8A",x"FE6A",x"FE8A",x"FE69",x"FE69",x"FE68",x"FE67",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE26",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE45",x"FE65",x"FE85",x"FE85",
									 x"E5A4",x"B404",x"6940",x"50A0",x"6120",x"6960",x"7160",x"7160",x"7180",x"79C2",
									 x"8B09",x"A490",x"BDD7",x"BE19",x"BDF8",x"BDF7",x"C617",x"C618",x"C639",x"C639",
									 x"C638",x"C638",x"D679",x"B596",x"944F",x"6AE8",x"4961",x"5160",x"59A0",x"59E0",
									 x"6A20",x"7241",x"8261",x"8261",x"8A81",x"9281",x"8A61",x"8A62",x"8A62",x"8240",
									 x"8AC0",x"9340",x"A440",x"D604",x"FF67",x"FFA6",x"FFA6",x"FF46",x"FF05",x"FEE5",
									 x"FEC5",x"FEA5",x"FEA5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE25",x"FE25",x"FE04",
									 x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD64",x"FD44",x"F503",x"FCE3",x"FCA3",x"F464",
									 x"E4A6",x"D50D",x"CD95",x"C5D7",x"BE17",x"CE7A",x"DEDB",x"EF3D",x"F79E",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F7FF",x"FFFF",x"FFDD",
									 x"FEF8",x"ED6F",x"F4A9",x"F403",x"F423",x"FC63",x"F483",x"FCC4",x"FCE4",x"FD04",
									 x"FD24",x"FD64",x"FD64",x"FD85",x"FD65",x"FDA4",x"FDC5",x"FDEA",x"FE6F",x"FED2",
									 x"FF35",x"FF57",x"FF57",x"FF56",x"FF56",x"FF36",x"FF36",x"FF35",x"FF35",x"FF15",
									 x"FF14",x"FF34",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FF11",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FE8C",x"FEAB",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",
									 x"FE69",x"FE68",x"FE68",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE46",x"FE26",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE65",x"FE65",x"FE85",x"EDC4",x"C464",x"71A0",x"58C0",
									 x"5900",x"6940",x"7160",x"7180",x"7160",x"7182",x"82C8",x"A46F",x"BDB6",x"C639",
									 x"BE19",x"BE18",x"C617",x"C618",x"C638",x"C618",x"C618",x"C638",x"CE79",x"C618",
									 x"AD53",x"83AC",x"4182",x"4960",x"51A0",x"59E0",x"6A20",x"7240",x"7A61",x"8281",
									 x"8A81",x"92A1",x"92A2",x"9282",x"9282",x"8A61",x"8261",x"8AC1",x"9B62",x"BCE5",
									 x"E686",x"F746",x"FF86",x"FF86",x"FF46",x"FF05",x"FEE5",x"FEC5",x"FEC5",x"FEC5",
									 x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",
									 x"FE65",x"FE65",x"FE65",x"FE45",x"FE25",x"FE05",x"FE04",x"FDE4",x"FDC4",x"FDA4",
									 x"FD84",x"FD64",x"FD24",x"FD04",x"FCC3",x"F482",x"EC84",x"E4A9",x"DD51",x"CDD5",
									 x"BDF5",x"C639",x"D69A",x"DEFB",x"EF7D",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF7B",x"F613",x"ECAA",x"F425",x"FC02",
									 x"FC42",x"FC83",x"F4C3",x"F4E3",x"FD04",x"FD24",x"FD44",x"FD64",x"FD84",x"FD85",
									 x"FD85",x"FDC5",x"F5E7",x"FE2E",x"FEB3",x"FF15",x"FF56",x"FF37",x"FF57",x"FF56",
									 x"FF56",x"FF36",x"FF36",x"FF35",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FECF",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAB",
									 x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE69",x"FE68",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE45",x"FE45",
									 x"FE65",x"FE85",x"EE04",x"CCC4",x"8260",x"6120",x"5900",x"6140",x"7160",x"7180",
									 x"7160",x"6961",x"7AA7",x"9C4E",x"BDD6",x"C639",x"BE18",x"BE17",x"C618",x"C618",
									 x"C638",x"C638",x"C638",x"C638",x"CE39",x"CE5A",x"CE59",x"9CD1",x"5205",x"4981",
									 x"4980",x"51C0",x"6200",x"6A40",x"7A61",x"8281",x"8AA1",x"92A1",x"92C1",x"9AC1",
									 x"9AC2",x"9AC2",x"92A1",x"8A81",x"8AA1",x"9B42",x"B483",x"DE05",x"F727",x"FF87",
									 x"FF67",x"FF46",x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE45",
									 x"FE45",x"FE25",x"FE05",x"FE04",x"FDC4",x"FDA4",x"FDA4",x"F584",x"FD64",x"FD24",
									 x"FCE3",x"F482",x"F463",x"EC87",x"E4ED",x"D592",x"BDB4",x"C618",x"CE79",x"D6BA",
									 x"EF5D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDD",x"FE96",x"ED0C",x"EC26",x"F3E3",x"F422",x"F483",x"F4C2",x"F4E3",x"FD04",
									 x"FD24",x"FD44",x"FD65",x"FD85",x"F584",x"F5A4",x"FDA6",x"FDE7",x"FE4B",x"FED2",
									 x"FF17",x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF35",
									 x"FF35",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAB",x"FE8B",x"FE8B",x"FE8B",x"FE8A",
									 x"FE6A",x"FE8A",x"FE89",x"FE68",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE45",x"FE45",x"FE65",x"FE85",x"F645",x"DD64",
									 x"9B21",x"6981",x"58E1",x"6100",x"6960",x"6960",x"6940",x"6121",x"7266",x"8BED",
									 x"B5B5",x"C638",x"BE18",x"BE18",x"C638",x"CE39",x"CE58",x"CE58",x"C638",x"C638",
									 x"C639",x"D69A",x"D6DB",x"B595",x"6AE9",x"51C2",x"4140",x"51A0",x"59E0",x"6A20",
									 x"7241",x"8281",x"8AA1",x"92A1",x"92C1",x"9AE1",x"A2E1",x"A2E1",x"A2E1",x"9AC1",
									 x"92A1",x"92A1",x"92E0",x"A401",x"BD02",x"E685",x"FF47",x"FF87",x"FF66",x"FF45",
									 x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",
									 x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",x"FE25",x"FE25",x"FE05",
									 x"FDE4",x"FDC4",x"FDC4",x"F584",x"FD84",x"FD44",x"FD03",x"FCC3",x"F483",x"F465",
									 x"E4A9",x"DD0E",x"CD72",x"BDF7",x"BDF7",x"CE59",x"DEFB",x"EF9E",x"FFBF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FF5B",x"F612",x"F4A8",x"F404",
									 x"F403",x"F463",x"F4A3",x"F4C2",x"F4E3",x"FD03",x"FD24",x"FD64",x"FD85",x"FD85",
									 x"F5A3",x"FDA4",x"FDC8",x"FE0A",x"FE8E",x"FF15",x"FF38",x"FF57",x"FF57",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF35",x"FF35",x"FF35",x"FF35",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FE8C",x"FEAB",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE6A",x"FE8A",x"FE89",x"FE68",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE45",x"FE45",x"FE65",x"FE65",x"FE65",x"EDC4",x"ABA2",x"71C2",x"58C0",x"58E0",
									 x"6940",x"6960",x"6961",x"6121",x"7246",x"83AB",x"AD74",x"BE18",x"BE18",x"C638",
									 x"C638",x"CE39",x"CE38",x"C638",x"CE59",x"CE59",x"C638",x"CE9A",x"D6DB",x"BDD7",
									 x"838C",x"59E4",x"4940",x"4960",x"59C0",x"6221",x"7221",x"7A61",x"8A81",x"92A1",
									 x"92C2",x"9AE2",x"A2E1",x"A2E0",x"A2E1",x"A302",x"9AE1",x"92A0",x"8A81",x"9301",
									 x"9BC1",x"CDA4",x"EEE6",x"FF88",x"FF87",x"FF66",x"FF25",x"FEE5",x"FEE5",x"FEE5",
									 x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",
									 x"FE85",x"FE65",x"FE45",x"FE45",x"FE25",x"FE05",x"FDE4",x"FDE5",x"FDC4",x"F5A4",
									 x"FD84",x"FD44",x"FD23",x"F4E3",x"F4C3",x"F4A3",x"ECA6",x"E4CA",x"DD30",x"BDD6",
									 x"BDD6",x"C638",x"D6BA",x"EF5D",x"FFBE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFBD",x"FED6",x"FD6D",x"F445",x"F403",x"F423",x"F463",x"F4C4",x"F4E3",
									 x"F503",x"F523",x"FD44",x"FD65",x"FD85",x"FD85",x"F584",x"FDA5",x"FE0A",x"FE8E",
									 x"FF12",x"FF56",x"FF58",x"FF57",x"FF57",x"FF56",x"FF36",x"FF56",x"FF36",x"FF36",
									 x"FF35",x"FF35",x"FF35",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF33",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAB",x"FE8B",x"FE8B",
									 x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE69",x"FE68",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"EE05",x"B402",x"7A01",x"58C0",x"58E0",x"7161",x"7161",x"6961",x"5920",
									 x"6A24",x"8349",x"AD12",x"C5F7",x"C618",x"C638",x"C638",x"C638",x"CE59",x"CE59",
									 x"CE59",x"CE59",x"CE59",x"CE79",x"D69A",x"CE59",x"9CB1",x"5205",x"4141",x"4960",
									 x"51A0",x"6201",x"6A21",x"7A61",x"8A81",x"92A1",x"92C2",x"9B02",x"A301",x"AB01",
									 x"AB01",x"A302",x"A302",x"A2E2",x"92A1",x"92C1",x"9300",x"AC02",x"CD64",x"E686",
									 x"F767",x"FFA7",x"FF66",x"FF26",x"FF06",x"FF05",x"FF05",x"FEE5",x"FEC5",x"FEE5",
									 x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",
									 x"FE45",x"FE25",x"FE04",x"FDE4",x"FDE4",x"FDA4",x"FDA4",x"FD84",x"FD43",x"FD03",
									 x"F4C3",x"F4A3",x"ECA4",x"ECA7",x"E4EC",x"CDB3",x"C5F7",x"C618",x"D678",x"E71B",
									 x"EF7E",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FEF8",x"F5D0",x"F4A8",
									 x"EC03",x"F423",x"F443",x"F483",x"FCC4",x"F4E4",x"F523",x"FD24",x"FD45",x"FD65",
									 x"FD84",x"FDA5",x"FD85",x"FDC8",x"FE6F",x"FEF3",x"FF56",x"FF78",x"FF57",x"FF57",
									 x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF35",x"FF35",x"FF35",x"FF35",x"FF35",
									 x"FF35",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",
									 x"FE8C",x"FE8C",x"FE8C",x"FEAB",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE69",
									 x"FE68",x"FE68",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE65",x"FE65",x"FE65",x"FEA6",x"F646",x"C4A4",x"8AA2",
									 x"58E0",x"50A0",x"6940",x"6960",x"6981",x"5940",x"61E3",x"7AC6",x"ACAF",x"BDB5",
									 x"C618",x"C639",x"CE38",x"C658",x"CE59",x"CE59",x"CE79",x"CE79",x"CE59",x"CE79",
									 x"CE7A",x"D6BB",x"BDF6",x"62E9",x"4182",x"4140",x"51A0",x"59E1",x"6221",x"7261",
									 x"8281",x"9281",x"92C1",x"9B02",x"A301",x"AB21",x"AB21",x"AB21",x"AB22",x"AB22",
									 x"A302",x"92E1",x"8AC0",x"9301",x"A3E1",x"BD03",x"DE65",x"F767",x"FF86",x"FF66",
									 x"FF26",x"FF25",x"FEE5",x"FEC5",x"FEC5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",
									 x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE05",x"FE04",
									 x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD63",x"FD24",x"FCE4",x"FCC3",x"F483",x"EC85",
									 x"E4A8",x"D550",x"CDD6",x"C5F8",x"C617",x"DEBA",x"E73D",x"F79E",x"FFDF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFDE",x"FF5B",x"FE74",x"F50C",x"F425",x"F423",x"F463",x"F463",x"F4A3",
									 x"FCE4",x"F504",x"FD24",x"FD45",x"FD65",x"FD64",x"FDA4",x"FDA5",x"FDC7",x"FE0C",
									 x"FED3",x"FF57",x"FF78",x"FF58",x"FF37",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF35",x"FF35",x"FF35",x"FF35",x"FF35",x"FF35",x"FF54",x"FF34",x"FF34",
									 x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FECF",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8C",x"FE8C",x"FE8C",x"FEAB",
									 x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE69",x"FE68",x"FE68",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE65",
									 x"FE65",x"FE65",x"FEA5",x"F685",x"CD24",x"9302",x"5920",x"50A0",x"6940",x"6960",
									 x"6980",x"5940",x"61C1",x"7265",x"A44E",x"BD94",x"C638",x"CE3A",x"CE59",x"CE58",
									 x"CE59",x"CE59",x"CE79",x"CE79",x"CE59",x"CE79",x"D69A",x"DEDB",x"C617",x"734B",
									 x"49E4",x"4140",x"4980",x"51C1",x"6200",x"7241",x"8261",x"8A81",x"92C1",x"9B01",
									 x"A301",x"AB22",x"AB42",x"AB22",x"AB42",x"AB42",x"AB42",x"A302",x"9AE1",x"92C0",
									 x"9300",x"9360",x"B503",x"E6C6",x"F767",x"FFA6",x"FF66",x"FF26",x"FF05",x"FEE5",
									 x"FEC5",x"FEE5",x"FEE6",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",
									 x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE25",x"FE04",x"FDE4",x"FDC4",x"FDA4",
									 x"FD64",x"FD44",x"FD04",x"FCE3",x"F4A2",x"F483",x"EC86",x"D4EC",x"CD93",x"BDD7",
									 x"BDF7",x"CE79",x"DEFB",x"EF5D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FEF8",x"FDF1",
									 x"F4A9",x"EC04",x"F422",x"F483",x"F483",x"F4C3",x"FD04",x"F504",x"F524",x"FD65",
									 x"FD65",x"FD64",x"FDA4",x"FDC6",x"FDE9",x"FE8F",x"FF15",x"FF79",x"FF78",x"FF57",
									 x"FF37",x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",x"FF36",x"FF35",x"FF35",x"FF35",
									 x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FE8C",x"FE8C",x"FE8C",x"FE8C",x"FEAB",x"FE8B",x"FE8B",x"FE8A",x"FE8A",
									 x"FE8A",x"FE69",x"FE68",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE65",x"FE65",x"FE65",x"FEC5",x"FEA5",
									 x"D564",x"9B62",x"6160",x"50C0",x"6120",x"6960",x"6980",x"6160",x"6180",x"6A03",
									 x"9C0D",x"B553",x"BE18",x"CE5A",x"CE59",x"CE59",x"CE59",x"CE79",x"CE79",x"CE79",
									 x"CE79",x"CE79",x"CE99",x"DEDB",x"CE58",x"83EE",x"5A66",x"3961",x"4160",x"51A1",
									 x"59E1",x"6A41",x"7A61",x"8A81",x"92C1",x"9B02",x"A301",x"AB21",x"AB42",x"AB42",
									 x"AB62",x"AB41",x"AB41",x"A321",x"A322",x"9AC1",x"92E1",x"9301",x"AC02",x"CDA5",
									 x"E6C6",x"F766",x"FF86",x"FF46",x"FF25",x"FF05",x"FEE5",x"FEE5",x"FEE6",x"FEE5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",
									 x"FE24",x"FE25",x"FE24",x"FDE4",x"FDE4",x"FDA4",x"FD84",x"FD64",x"FD24",x"FD03",
									 x"FCC2",x"FCA3",x"F485",x"DCC9",x"DD50",x"C595",x"BDD7",x"C658",x"D699",x"E71C",
									 x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FF7C",x"FE54",x"F50B",x"EC46",x"EC23",x"F462",x"F4A3",
									 x"F4A3",x"FCE3",x"FD24",x"FD44",x"FD44",x"FD65",x"FD65",x"FD84",x"FDC6",x"FE09",
									 x"FE4D",x"FEF2",x"FF57",x"FF79",x"FF58",x"FF56",x"FF36",x"FF57",x"FF57",x"FF57",
									 x"FF56",x"FF56",x"FF36",x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF55",x"FF54",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8C",x"FE8C",
									 x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE69",x"FE68",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE45",x"FE65",x"FE85",x"FEA5",x"FEC5",x"DDA4",x"ABE2",x"71E0",x"5900",
									 x"5900",x"6140",x"6960",x"6980",x"6180",x"69C2",x"93AC",x"B533",x"BE18",x"CE5A",
									 x"CE39",x"CE58",x"CE79",x"CE79",x"CE79",x"D69A",x"D69A",x"D69A",x"CE79",x"D6DA",
									 x"D69A",x"A4F2",x"7B6B",x"41A2",x"4140",x"49A1",x"59E1",x"6221",x"7261",x"8281",
									 x"92C1",x"9B02",x"A302",x"AB21",x"AB62",x"AB62",x"B362",x"AB61",x"AB61",x"AB41",
									 x"AB42",x"AB22",x"9B02",x"92E1",x"9321",x"A3E2",x"C544",x"E686",x"FF87",x"FFA7",
									 x"FF66",x"FF25",x"FF05",x"FEE5",x"FEE6",x"FEE5",x"FEE5",x"FEC5",x"FEC6",x"FEC5",
									 x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",x"FE45",x"FE25",x"FE04",
									 x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD44",x"FD23",x"FCE2",x"F4A2",x"F463",x"ECA6",
									 x"E4EB",x"D551",x"C5D6",x"BE17",x"C658",x"DEDB",x"EF5D",x"FFDF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"FED8",
									 x"F56E",x"EC46",x"F423",x"F441",x"F482",x"FCC3",x"F4C3",x"FD04",x"FD24",x"FD45",
									 x"FD65",x"FD85",x"FD85",x"FD85",x"FDE7",x"FE4C",x"FEB1",x"FF36",x"FF58",x"FF59",
									 x"FF38",x"FF37",x"FF37",x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",x"FF36",x"FF56",
									 x"FF56",x"FF56",x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8C",x"FE8C",x"FE8C",x"FE8B",x"FE8B",x"FE8B",
									 x"FE8A",x"FE8A",x"FE69",x"FE49",x"FE48",x"FE47",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE45",x"FE65",x"FE65",
									 x"FE86",x"FEA5",x"EE04",x"BC84",x"8A82",x"6120",x"50C0",x"6121",x"6960",x"6980",
									 x"6140",x"6182",x"934B",x"AD13",x"C638",x"CE7A",x"CE59",x"CE78",x"CE79",x"CE79",
									 x"D69A",x"D69A",x"D69A",x"D69A",x"CE99",x"D6BA",x"D6BA",x"C617",x"9C90",x"49E3",
									 x"3920",x"4981",x"51C0",x"6200",x"7261",x"7A81",x"8AA1",x"9AE2",x"A301",x"AB21",
									 x"AB62",x"B362",x"B382",x"B382",x"B382",x"B381",x"AB62",x"AB62",x"AB62",x"A322",
									 x"92E1",x"9300",x"A3E1",x"BCE3",x"E6C6",x"F786",x"FFA6",x"FF45",x"FF25",x"FF06",
									 x"FF06",x"FEE5",x"FEE5",x"FEE5",x"FEC6",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",
									 x"FE85",x"FE65",x"FE45",x"FE45",x"FE45",x"FE04",x"FE05",x"FDE4",x"FDC4",x"FDA4",
									 x"FD64",x"FD64",x"F503",x"F4E3",x"F484",x"EC85",x"EC88",x"DD0E",x"CDB4",x"B5F7",
									 x"BE38",x"CE79",x"E71C",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF5B",x"FE54",x"F4CA",x"EBE3",x"F422",x"F462",
									 x"FCA3",x"FCC3",x"FCE4",x"F504",x"FD24",x"FD45",x"FD65",x"FD85",x"FD84",x"FDC6",
									 x"FE2B",x"FEB0",x"FF15",x"FF58",x"FF58",x"FF58",x"FF58",x"FF58",x"FF37",x"FF57",
									 x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF55",
									 x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FE8C",x"FE8C",x"FE8C",x"FEAB",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE69",x"FE68",
									 x"FE67",x"FE47",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE66",x"FE46",x"FE46",x"FE65",x"FE65",x"FE65",x"FE86",x"FEA6",x"F645",x"CD03",
									 x"9302",x"6140",x"50A0",x"6121",x"6960",x"6960",x"5920",x"5962",x"8B2A",x"ACF3",
									 x"C638",x"CE9A",x"CE59",x"CE79",x"CE79",x"D69A",x"D69A",x"D69A",x"D69A",x"D69A",
									 x"D699",x"D6BA",x"D6BB",x"D6BA",x"AD53",x"5245",x"3120",x"4160",x"51A0",x"6201",
									 x"7261",x"7A81",x"8AA1",x"92E1",x"9AE1",x"AB21",x"B342",x"B362",x"B382",x"B382",
									 x"B3A2",x"B382",x"B382",x"AB62",x"AB62",x"AB62",x"A322",x"92E1",x"9321",x"9BC2",
									 x"CDA5",x"E6C5",x"FF87",x"FFA6",x"FF86",x"FF26",x"FF06",x"FEE5",x"FEE5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE45",
									 x"FE44",x"FE24",x"FE05",x"FE04",x"FDE4",x"FDC4",x"FDA4",x"FD64",x"FD24",x"FD04",
									 x"F4C4",x"EC83",x"F465",x"ECAB",x"D572",x"BDD6",x"B5F7",x"C638",x"D6DB",x"EF5D",
									 x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBD",
									 x"F6F9",x"F5D1",x"F467",x"F3E3",x"F423",x"F463",x"F483",x"FCC3",x"FD04",x"FD24",
									 x"FD24",x"FD44",x"FD65",x"FD85",x"FDA4",x"FDE7",x"FE6E",x"FEF3",x"FF57",x"FF58",
									 x"FF58",x"FF78",x"FF58",x"FF78",x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8C",x"FE8C",x"FEAB",
									 x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE69",x"FE68",x"FE67",x"FE47",x"FE67",x"FE67",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE65",
									 x"FE65",x"FE65",x"FEA5",x"FEA6",x"FE65",x"D543",x"A382",x"6160",x"50A0",x"6100",
									 x"6960",x"6960",x"5920",x"5942",x"832A",x"ACD1",x"C617",x"CE7A",x"CE7A",x"CE7A",
									 x"CE79",x"D69A",x"D69A",x"D69A",x"D69A",x"D6BA",x"D69A",x"D6BA",x"DEDC",x"E71C",
									 x"BDD5",x"62A7",x"3961",x"4160",x"51A0",x"61E1",x"7241",x"7260",x"82A1",x"92E1",
									 x"9B01",x"AB21",x"B342",x"B362",x"B382",x"BB82",x"BBA2",x"BBA2",x"B382",x"B382",
									 x"AB62",x"AB62",x"AB42",x"9B02",x"92C1",x"9301",x"AC43",x"D5C4",x"F747",x"FFE7",
									 x"FFC6",x"FF46",x"FF26",x"FF05",x"FF05",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE45",x"FE45",x"FE25",x"FE25",x"FE04",
									 x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD44",x"FD24",x"F4E3",x"F4A2",x"F463",x"ECA7",
									 x"D52E",x"C5B4",x"BDF7",x"BDF8",x"CE79",x"E73C",x"EF9E",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",x"FF5A",x"F634",x"ECEC",x"F425",x"F403",
									 x"F443",x"F483",x"F4A3",x"FCE4",x"FD04",x"FD44",x"FD44",x"FD65",x"FD65",x"FD85",
									 x"FDC6",x"FE2B",x"FEB1",x"FF36",x"FF78",x"FF78",x"FF58",x"FF78",x"FF57",x"FF57",
									 x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",
									 x"FF55",x"FF55",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FE8C",x"FE8C",x"FE8C",x"FEAB",x"FE8B",x"FE8B",x"FE8B",x"FE8A",
									 x"FE69",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE65",x"FE65",x"FE65",x"FE85",x"FEA6",
									 x"FEA6",x"DDA4",x"ABE3",x"6980",x"4880",x"5900",x"6960",x"6981",x"5920",x"5940",
									 x"7AE8",x"A46F",x"BDD6",x"CE7A",x"CE7A",x"CE7A",x"D69A",x"D69A",x"D6BA",x"D6BA",
									 x"D6BA",x"D6BA",x"D6BA",x"D6BB",x"DEDB",x"E71C",x"C5F6",x"734B",x"49C3",x"4161",
									 x"4980",x"59E0",x"6A41",x"7261",x"8281",x"92C2",x"9AE1",x"AB22",x"B342",x"B362",
									 x"B362",x"BB82",x"BBA2",x"BBA2",x"BBA2",x"B382",x"B382",x"B382",x"B383",x"AB43",
									 x"A322",x"92E1",x"9321",x"B463",x"CDE4",x"F746",x"FFC6",x"FFA6",x"FF66",x"FF26",
									 x"FF05",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",
									 x"FE65",x"FE65",x"FE65",x"FE45",x"FE25",x"FE04",x"FDE4",x"FDE4",x"FDC4",x"FD84",
									 x"FD64",x"FD44",x"FD03",x"F4E2",x"F4A2",x"ECA4",x"D4EA",x"CDB2",x"C5F7",x"BDD7",
									 x"C658",x"DEFB",x"E75C",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FF9C",x"FEB6",x"F58F",x"EC47",x"F403",x"F422",x"F463",x"F4A4",x"FCE4",x"FD04",
									 x"FD24",x"FD44",x"FD65",x"FD64",x"FD84",x"FDA5",x"FE09",x"FE6F",x"FF15",x"FF58",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF57",x"FF57",x"FF57",x"FF57",x"FF57",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FE8C",
									 x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE6A",x"FE69",x"FE68",x"FE47",x"FE47",
									 x"FE48",x"FE48",x"FE48",x"FE67",x"FE67",x"FE47",x"FE47",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE65",x"FE65",x"FE65",x"FE85",x"FE86",x"FEC6",x"E5E4",x"BC43",x"71C0",
									 x"4880",x"5900",x"6961",x"6981",x"6140",x"5940",x"7A85",x"9C0D",x"BD95",x"CE79",
									 x"CE9A",x"CE7A",x"D69A",x"D69A",x"D6BA",x"D6BA",x"D6BA",x"D6BA",x"D69A",x"DEDB",
									 x"DEDB",x"E71C",x"CE58",x"946F",x"5245",x"3941",x"4960",x"59C0",x"6A41",x"6A40",
									 x"7A81",x"8AC2",x"9AE1",x"A321",x"AB42",x"B362",x"B362",x"BB82",x"BBA2",x"BBA2",
									 x"BBA2",x"BBA2",x"B3A2",x"B382",x"B382",x"AB42",x"AB42",x"9B22",x"92C1",x"9B42",
									 x"B482",x"DE65",x"FF86",x"FFA7",x"FF86",x"FF46",x"FF25",x"FEE5",x"FEE5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",
									 x"FE45",x"FE25",x"FE04",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD64",x"FD23",x"FCE3",
									 x"F4A2",x"EC83",x"DCC7",x"D56F",x"C5B6",x"BDB6",x"C638",x"D6BA",x"DF1B",x"F79E",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF7B",x"FE33",x"F50B",x"EC25",
									 x"F402",x"F442",x"F483",x"F4A3",x"FCE4",x"FD24",x"FD24",x"FD64",x"FD84",x"FD84",
									 x"FD85",x"FDC7",x"FE4C",x"FED3",x"FF38",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAB",x"FEAB",x"FEAB",
									 x"FE8B",x"FE8A",x"FE89",x"FE68",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE67",
									 x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FEA6",x"FEC6",x"E624",x"C4A3",x"8240",x"48A0",x"5900",x"6140",x"6960",
									 x"6140",x"6160",x"7243",x"93AB",x"B553",x"C638",x"CE9A",x"CE9A",x"D69A",x"D69A",
									 x"D6BA",x"D6BA",x"D6BA",x"D6BA",x"DEDA",x"DEDB",x"DEBB",x"E6FC",x"D699",x"AD54",
									 x"62C8",x"3941",x"4140",x"51A0",x"6200",x"6A40",x"7A61",x"8AC2",x"9AE1",x"A301",
									 x"AB42",x"B362",x"BB62",x"BB82",x"BBA2",x"BBA2",x"BBA2",x"BBA2",x"BBC3",x"B3A2",
									 x"B382",x"B382",x"AB62",x"AB62",x"9AE2",x"9B02",x"9BA1",x"C544",x"EEC6",x"F767",
									 x"FF87",x"FF45",x"FF46",x"FF05",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",x"FE25",x"FE04",x"FE04",
									 x"FDE4",x"FDC4",x"FD84",x"FD64",x"FD43",x"F503",x"F4A3",x"F483",x"EC85",x"DD0D",
									 x"CD74",x"C5B6",x"C617",x"CE79",x"D6DA",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFDF",x"FF19",x"F58F",x"EC88",x"EC24",x"F422",x"F463",x"F4A3",x"FCC3",
									 x"FCE3",x"FD24",x"FD44",x"FD64",x"FDA5",x"FD84",x"FD86",x"FE09",x"FEAF",x"FF15",
									 x"FF5A",x"FF59",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",
									 x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF55",
									 x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FECC",x"FECB",x"FECB",x"FEAB",
									 x"FEAB",x"FEAB",x"FEAB",x"FECB",x"FECC",x"FECC",x"FECB",x"FECA",x"FEA9",x"FEA8",
									 x"FEA8",x"FEA8",x"FEA8",x"FE88",x"FE87",x"FE87",x"FE67",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FEA6",x"FEC6",x"EE44",
									 x"D524",x"8AA1",x"50E0",x"5900",x"6120",x"6960",x"6160",x"6160",x"7201",x"8B48",
									 x"ACF1",x"C617",x"CE9A",x"CE9A",x"D69A",x"D6BA",x"D6BA",x"D6BA",x"D6BA",x"D6BA",
									 x"DEDA",x"D6BB",x"DEBB",x"DEFC",x"DEDB",x"CE59",x"7B6B",x"3941",x"4120",x"51A0",
									 x"6200",x"6A40",x"7A61",x"8AC2",x"92C1",x"A301",x"AB42",x"B362",x"BB82",x"BB82",
									 x"C3A2",x"C3C2",x"BBC2",x"BBC2",x"BBC3",x"B3C3",x"B3A2",x"B382",x"B382",x"ABA2",
									 x"A322",x"9B02",x"9321",x"A422",x"CDA5",x"EEE6",x"FFA7",x"FF86",x"FF46",x"FF25",
									 x"FF05",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",
									 x"FE85",x"FE65",x"FE45",x"FE45",x"FE24",x"FE05",x"FDE4",x"FDC4",x"FDA4",x"FD84",
									 x"FD43",x"FD03",x"F4C3",x"F483",x"F464",x"DCC9",x"CD51",x"C5B6",x"BDD6",x"C638",
									 x"CE9A",x"E73C",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"F79D",x"FE95",x"ECAA",
									 x"EC25",x"EC23",x"F443",x"F483",x"F4A3",x"FCC3",x"FD03",x"FD44",x"F544",x"FD64",
									 x"FDA5",x"FDA5",x"FDC7",x"FE4C",x"FEF3",x"FF58",x"FF7A",x"FF79",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FEAD",x"FEAD",
									 x"FEAD",x"FE8C",x"FEAD",x"FEAC",x"FECC",x"FECB",x"FEAB",x"F68B",x"F66C",x"EE6B",
									 x"EE6B",x"EE6B",x"F66B",x"EE6A",x"EE6A",x"EE68",x"F688",x"F688",x"F6A8",x"FEA9",
									 x"FEA8",x"FEA8",x"FEA8",x"FE87",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE85",x"FEC6",x"EE64",x"DD64",x"9B01",x"5940",x"5900",
									 x"5900",x"6940",x"6160",x"6160",x"69C1",x"82E7",x"ACB0",x"C5F7",x"D69B",x"CE9A",
									 x"D69A",x"D6BA",x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"D6BA",x"D6BA",x"DEDB",x"DEDB",
									 x"E71C",x"E71C",x"8C2E",x"4182",x"4140",x"51A0",x"59E0",x"6220",x"7261",x"82C2",
									 x"92E1",x"9B01",x"AB41",x"B362",x"B362",x"BB82",x"C3C2",x"C3C2",x"C3C2",x"BBC2",
									 x"BBE3",x"BBC3",x"BBC2",x"B3A2",x"B3A2",x"ABA2",x"AB62",x"A362",x"9301",x"9341",
									 x"AC43",x"CDC4",x"EF06",x"FFA6",x"FF65",x"FF46",x"FF05",x"FEE5",x"FEE5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",
									 x"FE25",x"FE05",x"FDE4",x"FDE4",x"FDA4",x"FDA4",x"FD63",x"FD23",x"F4E3",x"F4C3",
									 x"EC83",x"E4A7",x"DD0D",x"CD94",x"BDB5",x"BE17",x"C679",x"DEFB",x"F77E",x"F7BF",
									 x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFBE",x"FF3A",x"F632",x"EC47",x"F403",x"F423",x"F463",x"F4A3",
									 x"F4C3",x"F4E3",x"FD24",x"FD45",x"F565",x"FD65",x"FDA5",x"FDC6",x"FDE9",x"FE8F",
									 x"FF36",x"FF79",x"FF79",x"FF79",x"FF78",x"FF58",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",
									 x"FF55",x"FF55",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FECD",x"FEAD",
									 x"FECD",x"FEAC",x"EE4B",x"DDAA",x"CD29",x"BCE7",x"B486",x"B466",x"AC25",x"A404",
									 x"A404",x"AC44",x"BCC5",x"C526",x"D586",x"E628",x"F6A9",x"FEEA",x"FF09",x"FEC8",
									 x"FEA8",x"FE88",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",
									 x"FEA6",x"F684",x"E5C4",x"A362",x"6180",x"5900",x"5900",x"6140",x"6960",x"6140",
									 x"6181",x"7A85",x"A46F",x"C5F8",x"D69B",x"D6BA",x"D69A",x"D6BA",x"DEDB",x"DEDB",
									 x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"E71C",x"E73C",x"9490",x"4A04",
									 x"4181",x"4980",x"59E0",x"6200",x"7261",x"82C2",x"8AC1",x"9B01",x"A341",x"AB62",
									 x"B362",x"BB82",x"C3A2",x"C3C2",x"C3C2",x"C3E2",x"BBE2",x"BBE2",x"BBC2",x"BBC2",
									 x"B3C2",x"B3A2",x"AB82",x"AB62",x"9B41",x"9301",x"9B82",x"BCC4",x"DE45",x"FFA7",
									 x"FFA6",x"FF86",x"FF26",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",
									 x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE65",x"FE45",x"FE45",x"FE05",x"FE05",x"FDE4",
									 x"FDC4",x"FDA4",x"F584",x"FD44",x"F503",x"F4E3",x"ECA3",x"E486",x"E4AA",x"D550",
									 x"BD94",x"B5F7",x"C638",x"D69A",x"EF5D",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF9D",x"F6B7",
									 x"F58E",x"EC25",x"F403",x"F443",x"F483",x"F4A3",x"F4E4",x"FD04",x"FD24",x"FD65",
									 x"FD65",x"FD65",x"FD85",x"FDC7",x"FE2C",x"FEF2",x"FF98",x"FF99",x"FF79",x"FF78",
									 x"FF78",x"FF58",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",
									 x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FECC",x"FEAC",x"EE4C",x"DDCB",x"CD0A",x"B468",
									 x"9BC5",x"8B03",x"7AA2",x"7241",x"6A20",x"6A00",x"6A00",x"7261",x"8B02",x"9BA4",
									 x"AC45",x"CD27",x"E5E9",x"EE4A",x"F6CA",x"FF09",x"FF08",x"FEE8",x"FEA8",x"FE88",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FEA6",x"F684",x"EE04",x"ABC3",
									 x"71E0",x"5900",x"58E0",x"6140",x"6980",x"6140",x"6140",x"7245",x"9C4F",x"C5D7",
									 x"D6BB",x"D6DA",x"D69A",x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"DEDB",
									 x"DEDB",x"DEFB",x"E73C",x"E73C",x"A4D1",x"5A87",x"4182",x"4980",x"59E1",x"6220",
									 x"7261",x"82C2",x"8AC1",x"9301",x"A341",x"AB42",x"B362",x"BB82",x"BBA2",x"C3C2",
									 x"C3C2",x"C3E2",x"C3E2",x"BBE2",x"BBE2",x"BBC2",x"BBC2",x"B3C2",x"B3A2",x"AB82",
									 x"AB62",x"9B02",x"9322",x"AC02",x"C563",x"F746",x"FFC6",x"FFC7",x"FF46",x"FF05",
									 x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",
									 x"FE65",x"FE45",x"FE45",x"FE25",x"FE05",x"FDE5",x"FDC4",x"FDC4",x"FD84",x"FD64",
									 x"FD04",x"FCE3",x"F4A3",x"EC85",x"EC88",x"D50D",x"C593",x"BDF7",x"BDF8",x"CE79",
									 x"E71C",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF5B",x"F633",x"ECCA",x"EC03",x"EC02",x"F443",
									 x"F483",x"FCC4",x"FCE4",x"FD04",x"FD45",x"FD65",x"FD65",x"FD65",x"FD86",x"FDC9",
									 x"FE8F",x"FF55",x"FF99",x"FF99",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FEAC",x"FECD",x"FECD",
									 x"F66B",x"DDCA",x"B487",x"8B23",x"7242",x"7221",x"6A20",x"6A21",x"7201",x"7221",
									 x"7221",x"7221",x"7221",x"7241",x"7A61",x"7A81",x"7A81",x"82A1",x"8B01",x"9BA3",
									 x"C526",x"EE89",x"FF2A",x"FF49",x"FF29",x"FEC9",x"FE87",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE46",x"FE46",x"FE66",x"FE66",x"FE46",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE84",x"FEA6",x"FE84",x"F645",x"BC23",x"7A21",x"5920",x"50C0",x"6160",
									 x"6980",x"6140",x"5920",x"6A24",x"9C0E",x"C5D7",x"D6BB",x"D6BA",x"D6BA",x"DEDB",
									 x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"DEFB",x"E73C",x"E73C",
									 x"B574",x"734B",x"49E4",x"4140",x"51C0",x"5A00",x"6A41",x"7AA2",x"82C1",x"9301",
									 x"A322",x"AB42",x"B362",x"B3A2",x"BBC2",x"C3C2",x"C3C2",x"C3E2",x"C3E2",x"C3E2",
									 x"C3E2",x"BBE2",x"BBC2",x"BBC2",x"B3A2",x"B382",x"AB82",x"A343",x"9B22",x"9301",
									 x"AC41",x"D665",x"F786",x"FFE7",x"FF86",x"FF26",x"FF05",x"FF05",x"FEC5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",x"FE25",
									 x"FE25",x"FE05",x"FDE4",x"FDC4",x"FDA4",x"FD64",x"FD24",x"FD04",x"FCC3",x"F484",
									 x"F486",x"DCCA",x"CD71",x"C5D6",x"BDD7",x"C638",x"DEFB",x"EF5D",x"F7BE",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",
									 x"FEF8",x"F590",x"F467",x"EC23",x"F422",x"F463",x"FCA3",x"FCE4",x"FD04",x"FD24",
									 x"FD65",x"FD85",x"FD85",x"FD85",x"FDA7",x"F60B",x"FED2",x"FF77",x"FF99",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF57",x"FF57",x"FF56",x"FF56",x"FF36",x"FF36",x"FF36",x"FF55",x"FF55",x"FF55",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FF11",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECE",x"FECD",x"FEAD",x"FEAD",x"EE2C",x"C4E8",x"AC26",x"8B03",x"61E0",
									 x"5980",x"61C0",x"6A00",x"7221",x"7A41",x"7A61",x"8281",x"8281",x"8282",x"8281",
									 x"8281",x"8281",x"7A41",x"7200",x"7221",x"7A81",x"9383",x"C507",x"E649",x"EEEA",
									 x"FF4B",x"FF09",x"FEC8",x"FEA8",x"FE87",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE66",x"FE66",
									 x"FE46",x"FE46",x"FE46",x"FE65",x"FE65",x"FE65",x"FE64",x"FE64",x"FE86",x"FEA4",
									 x"F685",x"C483",x"8261",x"5940",x"50C0",x"6160",x"6980",x"6941",x"5900",x"6A04",
									 x"940D",x"C5B6",x"D6DB",x"D6BA",x"D6BA",x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"DEFB",
									 x"DEFB",x"DEFB",x"DEFB",x"E71C",x"E73C",x"E73C",x"BDD6",x"8C0E",x"5A26",x"3920",
									 x"51A0",x"59E0",x"6A41",x"7AA2",x"82C1",x"92E1",x"A322",x"AB42",x"AB62",x"B3A2",
									 x"BBA2",x"C3C2",x"C3C2",x"C3E2",x"C3E2",x"C3E2",x"C3E2",x"C3E2",x"BBE2",x"BBE3",
									 x"BBA2",x"B3A2",x"B3A2",x"AB83",x"A343",x"92E1",x"9B81",x"C544",x"E6E6",x"FFA7",
									 x"FF87",x"FF46",x"FF26",x"FF05",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FE85",x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE25",x"FDE4",x"FDE4",
									 x"FDC4",x"FD84",x"FD44",x"FD24",x"FCE3",x"F4A3",x"F464",x"E4A8",x"D54F",x"C5B5",
									 x"BDB6",x"C618",x"D6BA",x"E73C",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF7C",x"F655",x"F50C",x"F426",x"EC22",
									 x"F442",x"FC83",x"FCA3",x"FCE4",x"FD04",x"FD24",x"FD64",x"FD85",x"FD84",x"FDA5",
									 x"FDE9",x"FE6E",x"FF14",x"FF98",x"FF7A",x"FF79",x"FF78",x"FF58",x"FF78",x"FF58",
									 x"FF58",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",x"FF56",x"FF56",
									 x"FF36",x"FF36",x"FF36",x"FF55",x"FF55",x"FF55",x"FF35",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FEF2",x"FEF1",x"FEF1",x"FF11",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FEED",x"FECE",
									 x"EE4D",x"C50A",x"8B24",x"6A21",x"61E0",x"61E0",x"6A01",x"7221",x"7A41",x"7A61",
									 x"8281",x"82A1",x"8AA1",x"8AA1",x"8AA2",x"8AA2",x"8AA1",x"8AA1",x"8A82",x"8261",
									 x"8261",x"7A61",x"7240",x"9343",x"BCC6",x"D5E8",x"FF2B",x"FF4A",x"FF29",x"FEE8",
									 x"FEA8",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE64",x"FE66",x"FEA4",x"FEA5",x"CD04",x"8AA1",x"5940",
									 x"48A0",x"6140",x"6981",x"6941",x"58E0",x"61E4",x"93ED",x"BDB6",x"D6DB",x"D6BB",
									 x"D6BA",x"DEDB",x"DEFB",x"DEFB",x"DEDB",x"DEFB",x"DEFB",x"DEFB",x"E71C",x"E71C",
									 x"E73C",x"E73C",x"CE78",x"A512",x"6288",x"3100",x"4980",x"51E0",x"6A21",x"7A82",
									 x"82A1",x"92E1",x"A322",x"AB42",x"AB62",x"B3A2",x"BBC2",x"C3C2",x"C3C2",x"C3E2",
									 x"C3E2",x"C3E2",x"C3E2",x"C3E2",x"C3E2",x"BBE3",x"BBC2",x"B3C2",x"B3C2",x"ABA2",
									 x"A363",x"9B22",x"9B42",x"B443",x"DE25",x"EF26",x"FF87",x"FF86",x"FF46",x"FF05",
									 x"FF05",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",
									 x"FE65",x"FE45",x"FE45",x"FE25",x"FE04",x"FDE4",x"FDC4",x"FD83",x"FD64",x"FD24",
									 x"F4E3",x"F4A3",x"F484",x"EC87",x"D50D",x"C5B3",x"BDD5",x"C5F8",x"CE7A",x"DEFB",
									 x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FF3A",x"F5F1",x"F4A9",x"EC24",x"EC42",x"F462",x"F4A3",x"FCC4",x"FCE4",
									 x"FD04",x"FD24",x"FD64",x"FD85",x"FD84",x"FDC6",x"FE4C",x"FEB2",x"FF37",x"FF99",
									 x"FF79",x"FF79",x"FF78",x"FF58",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF55",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FF11",
									 x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FEAE",x"FEEE",x"FECD",x"EE4C",x"C4E9",x"8B05",x"61C1",x"5980",
									 x"61A0",x"6A00",x"7A41",x"7A81",x"8282",x"82A1",x"8AA1",x"8AC1",x"8AE1",x"92E1",
									 x"92E2",x"92C2",x"92C2",x"92C2",x"92C2",x"92E2",x"8AC1",x"8AA1",x"7A40",x"7A41",
									 x"8AE2",x"A403",x"DE29",x"FF6B",x"FF8B",x"FF29",x"FEC8",x"FE88",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FEA5",x"FEC5",x"D544",x"92E1",x"6161",x"48A0",x"6140",x"6980",x"6941",
									 x"5901",x"61C4",x"93AC",x"B594",x"D6DA",x"D6BB",x"D6BA",x"DEDB",x"DEFB",x"DEFB",
									 x"DEFB",x"DEFB",x"DEFB",x"DEFB",x"DEFB",x"E71C",x"E71C",x"E73C",x"DEDB",x"C5D6",
									 x"6AC9",x"30E0",x"4980",x"59E0",x"6220",x"7281",x"7AA1",x"8AE1",x"9B22",x"A342",
									 x"AB61",x"B3A2",x"BBA2",x"BBC2",x"C3C2",x"C3E2",x"C3E2",x"C3E2",x"C3E2",x"C3E2",
									 x"C3E2",x"C3E2",x"BBC2",x"BBE2",x"B3E2",x"B3C2",x"ABA2",x"A362",x"9301",x"A382",
									 x"C544",x"DE64",x"F767",x"FFA7",x"FF66",x"FF26",x"FF05",x"FEE5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",x"FE25",
									 x"FE04",x"FE04",x"FDE4",x"FDA3",x"FD84",x"FD44",x"F503",x"F4C3",x"F483",x"EC65",
									 x"DCCA",x"CD70",x"C5D5",x"BDF7",x"C639",x"DEBA",x"E73C",x"F7BE",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FED7",x"F54D",x"EC67",
									 x"EC43",x"EC42",x"F462",x"F4A3",x"FCC4",x"FD04",x"FD24",x"FD44",x"FD85",x"FD85",
									 x"FD85",x"FDC7",x"FE8E",x"FF15",x"FF79",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",
									 x"FF58",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF55",x"FF35",x"FF54",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FED0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FEEF",
									 x"EE4C",x"BCE8",x"9386",x"61A1",x"5180",x"61E0",x"7201",x"7A62",x"8282",x"8281",
									 x"8AA1",x"8AC1",x"92E1",x"92E1",x"92E1",x"9301",x"9B01",x"9AE2",x"9AE2",x"9AE2",
									 x"92E2",x"9B02",x"92E1",x"92E1",x"92C2",x"8241",x"79E0",x"7A80",x"AC84",x"E6AA",
									 x"FF8C",x"FF8A",x"FF09",x"FEA9",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE66",x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE66",x"FE85",x"FEC5",x"FEC6",x"D583",
									 x"9B41",x"6181",x"48A0",x"5940",x"6980",x"6961",x"5900",x"61A3",x"8B6A",x"AD52",
									 x"CEB9",x"D6BA",x"DEDA",x"DEDB",x"DEFB",x"DEFB",x"DEFB",x"DEFB",x"DEFB",x"DEFB",
									 x"DEFB",x"DEFB",x"E71C",x"E73C",x"E73C",x"D658",x"7B2B",x"3900",x"4960",x"51C0",
									 x"6200",x"7261",x"7AA1",x"8AC1",x"9B21",x"A341",x"AB61",x"B382",x"BBA1",x"BBC2",
									 x"C3C2",x"C3E2",x"C3E3",x"C3E3",x"C3E3",x"C3E3",x"C403",x"C3E2",x"BBE2",x"BBE2",
									 x"BBE2",x"B3C2",x"B3A2",x"ABA2",x"9B41",x"9321",x"AC22",x"C583",x"EF07",x"FFC7",
									 x"FFA6",x"FF66",x"FF05",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",
									 x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",x"FE24",x"FE04",x"FDE4",x"FDA4",
									 x"FD84",x"FD64",x"FD24",x"F4E3",x"F4A3",x"F464",x"E4A8",x"D52E",x"CDB4",x"BDD7",
									 x"C618",x"D67A",x"E6FC",x"F79E",x"F7DF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFE",x"FF9D",x"FE55",x"ECCA",x"EC45",x"EC23",x"F462",x"F483",x"FCA3",
									 x"FCE4",x"FD04",x"FD44",x"FD44",x"FD85",x"FD85",x"FD85",x"FDE9",x"FED1",x"FF57",
									 x"FF99",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF58",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF55",x"FF55",x"FF55",x"FF34",x"FF54",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FEEE",x"FECE",x"FEEE",x"DDCB",x"93A5",x"7284",x"5981",
									 x"61C0",x"6A20",x"7241",x"7A81",x"8281",x"82A1",x"8AC1",x"8AC1",x"92E1",x"92E1",
									 x"9B01",x"9B02",x"9B02",x"9B02",x"9B02",x"9B02",x"9B22",x"9B02",x"9B02",x"9B01",
									 x"9AE2",x"9282",x"8A41",x"8260",x"9342",x"CDA9",x"EF2B",x"FF8B",x"FF49",x"FEE9",
									 x"FE88",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE85",x"FEC5",x"FEC6",x"DDC4",x"A382",x"69A0",x"50C0",x"5920",
									 x"6960",x"6961",x"5920",x"69A2",x"8B49",x"AD11",x"CE99",x"D6BB",x"DEDB",x"DEFB",
									 x"DEFB",x"DEFB",x"DEFB",x"DEFB",x"E71C",x"E71C",x"E71C",x"E71C",x"E71C",x"E73C",
									 x"EF5D",x"DEBA",x"838C",x"3941",x"4960",x"51A0",x"5A00",x"6A61",x"7A81",x"8AC1",
									 x"9B21",x"A321",x"AB41",x"B382",x"BBA2",x"BBC2",x"C3C2",x"C3E2",x"C3E3",x"C3E3",
									 x"C3E3",x"C403",x"C403",x"C402",x"BBE2",x"BC02",x"BBE2",x"B3E2",x"B3C2",x"ABA2",
									 x"A361",x"9B41",x"9B82",x"AC83",x"DE66",x"FFA7",x"FFC6",x"FF86",x"FF25",x"FF05",
									 x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",
									 x"FE65",x"FE45",x"FE25",x"FE24",x"FE04",x"FDC4",x"FDA4",x"F584",x"FD44",x"FD03",
									 x"FCA3",x"F483",x"ECA7",x"DD0C",x"D5B3",x"C5D6",x"BE18",x"CE59",x"DEDB",x"EF7D",
									 x"F7DE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FF3B",x"F5D2",
									 x"EC48",x"F424",x"EC22",x"F462",x"F4A3",x"FCC3",x"FCE4",x"FD04",x"FD44",x"FD64",
									 x"FD65",x"FD85",x"F5A6",x"FE4C",x"FF14",x"FF98",x"FF99",x"FF79",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF35",
									 x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FEEF",x"FEEE",
									 x"FECE",x"F68D",x"BCE9",x"6A22",x"5981",x"59C1",x"6A00",x"7240",x"7A61",x"8281",
									 x"82A1",x"8AC1",x"8AC1",x"92E1",x"9301",x"9B01",x"9B02",x"9B22",x"A322",x"A322",
									 x"A322",x"A322",x"A322",x"9B02",x"9B02",x"9B01",x"9AE1",x"9AC2",x"92A2",x"8241",
									 x"8261",x"B486",x"D649",x"F76B",x"FFAB",x"FF2A",x"FEC8",x"FE67",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FEC5",
									 x"FEE6",x"E604",x"ABE2",x"7200",x"5100",x"5920",x"6160",x"6961",x"5900",x"6182",
									 x"8307",x"A4CF",x"CE78",x"D6BB",x"DEDB",x"DEFB",x"DEFB",x"E71C",x"E71C",x"E71C",
									 x"E71C",x"E71C",x"E71C",x"E71C",x"E71C",x"E73C",x"EF7D",x"DEDA",x"8BEE",x"4183",
									 x"4160",x"5180",x"59E0",x"6A61",x"7281",x"82C1",x"9301",x"A341",x"AB42",x"B382",
									 x"BBA2",x"BBC2",x"C3C2",x"C3E2",x"C3E3",x"C403",x"C403",x"C403",x"C402",x"C3E2",
									 x"BBE2",x"BC02",x"BC02",x"BBE2",x"BBE2",x"B3C2",x"B3A2",x"A341",x"9301",x"9BA2",
									 x"CD85",x"F747",x"FFC6",x"FFA6",x"FF45",x"FF05",x"FEE6",x"FEC6",x"FEC6",x"FEC5",
									 x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE25",
									 x"FE04",x"FDE4",x"F5C4",x"FDA4",x"FD64",x"FD03",x"FCC3",x"FC83",x"EC85",x"E4EA",
									 x"D550",x"C5B5",x"B5D7",x"C638",x"D6BA",x"EF5D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFE",x"FFBD",x"FEB8",x"F54E",x"EC26",x"F423",x"F442",x"F482",
									 x"F4A3",x"F4C3",x"FD04",x"FD24",x"FD64",x"FD85",x"FD85",x"FDA5",x"F5E7",x"FE8F",
									 x"FF37",x"FF79",x"FF99",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",
									 x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FF12",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FECF",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FEEE",x"FECE",x"E60C",x"A3E7",x"5181",
									 x"4900",x"61E1",x"7241",x"7A41",x"7A81",x"82A1",x"8AC1",x"8AE1",x"92E1",x"9301",
									 x"9B02",x"9B22",x"A322",x"A322",x"A322",x"A322",x"A322",x"A322",x"A322",x"A342",
									 x"A322",x"A321",x"9B01",x"9AE2",x"9AE2",x"8A81",x"8261",x"9BA4",x"B506",x"E6EA",
									 x"FFCB",x"FF4A",x"FEE9",x"FE87",x"FE47",x"FE47",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FEA4",x"FEE6",x"EE25",x"B443",x"8261",
									 x"5940",x"5900",x"6140",x"6960",x"5920",x"6981",x"7AA5",x"9C6C",x"C636",x"D6BB",
									 x"DEFB",x"DEFB",x"DEFB",x"E71C",x"E71C",x"E73C",x"E71C",x"E73C",x"E73C",x"E73C",
									 x"E73C",x"E73C",x"EF7D",x"DEFB",x"9490",x"4A05",x"4140",x"4960",x"59E0",x"6A41",
									 x"7261",x"82A1",x"9301",x"A342",x"AB42",x"B362",x"B3A2",x"BBC2",x"C3C2",x"C3E2",
									 x"C3E2",x"C402",x"CC03",x"C402",x"C402",x"C3E2",x"C402",x"C402",x"BC02",x"BBE2",
									 x"BBE2",x"B3E2",x"B3C2",x"AB62",x"9B02",x"9322",x"B483",x"DE66",x"F766",x"FFC6",
									 x"FF66",x"FF26",x"FF06",x"FEE6",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",x"FE04",x"FDE5",x"F5C4",x"FDA4",
									 x"FD64",x"FD23",x"FCE3",x"FCA3",x"F484",x"E4C8",x"DD2E",x"C593",x"BDD7",x"C638",
									 x"CE79",x"E73C",x"F77E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",x"F75C",
									 x"FE55",x"ECEC",x"EC04",x"F422",x"F462",x"F4A3",x"F4C3",x"F4E3",x"FD24",x"FD44",
									 x"FD64",x"FD85",x"FD85",x"F5A5",x"F628",x"FED1",x"FF39",x"FF7A",x"FF79",x"FF79",
									 x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",
									 x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECF",
									 x"FEEF",x"FECE",x"F68C",x"D54A",x"8B25",x"5181",x"4960",x"6200",x"7242",x"7A61",
									 x"82A1",x"82A1",x"8AE2",x"9301",x"9301",x"9B21",x"A322",x"A322",x"A322",x"A342",
									 x"A322",x"A342",x"A342",x"A342",x"A342",x"AB42",x"A342",x"A322",x"9B22",x"9B02",
									 x"9B02",x"92C1",x"8A80",x"8AE2",x"9BC3",x"DEAA",x"FFCC",x"FF8B",x"FF09",x"FE87",
									 x"FE67",x"FE47",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",
									 x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE85",x"FEA4",x"FEE6",x"EE45",x"C4A3",x"8AE1",x"6160",x"5900",x"6120",x"6960",
									 x"6140",x"6180",x"7263",x"940A",x"C616",x"D6BB",x"DEFB",x"DEFB",x"E71C",x"E73C",
									 x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"EF7D",x"DEFB",
									 x"A512",x"5A67",x"3940",x"4960",x"59E0",x"6A41",x"7261",x"82A1",x"92E1",x"9B21",
									 x"A322",x"AB62",x"B382",x"BBC2",x"C3C2",x"C3E2",x"C3E2",x"C402",x"CC02",x"C402",
									 x"C402",x"C402",x"C402",x"C403",x"C402",x"BC02",x"BBE2",x"BBE2",x"B3E2",x"ABA2",
									 x"A362",x"9B21",x"9BA0",x"CD84",x"EF06",x"FFA6",x"FF87",x"FF46",x"FF06",x"FEE5",
									 x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",
									 x"FE65",x"FE45",x"FE24",x"FDE5",x"FDE4",x"FDC4",x"FD84",x"F543",x"F503",x"F4C3",
									 x"F484",x"ECA7",x"DCEC",x"CD72",x"BDD6",x"BE18",x"C638",x"E6FB",x"EF5D",x"FFBF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FF3A",x"FDF1",x"ECA9",x"EC03",x"F422",
									 x"F462",x"F4A3",x"F4C3",x"F4E3",x"FD24",x"FD44",x"FD65",x"FD65",x"FD85",x"F5C6",
									 x"F62B",x"FEF4",x"FF5A",x"FF7A",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FEEF",x"FEEF",x"FECE",x"F68D",x"C4E9",
									 x"7AA3",x"5180",x"5180",x"6A20",x"7241",x"7A61",x"8281",x"8AA1",x"92E1",x"9302",
									 x"9B02",x"9B22",x"A322",x"A322",x"A342",x"AB42",x"AB42",x"AB42",x"AB42",x"AB42",
									 x"AB42",x"AB42",x"A342",x"A322",x"A322",x"9B01",x"9B01",x"92E1",x"8AA1",x"82A1",
									 x"8B21",x"DE69",x"FFCC",x"FF8B",x"FF09",x"FE88",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FEA5",x"FEC6",x"F665",
									 x"CCE4",x"9321",x"6980",x"5900",x"5920",x"6160",x"6140",x"6160",x"7222",x"93EA",
									 x"C615",x"D6BB",x"DEFB",x"E71C",x"E71C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",
									 x"E73C",x"E73C",x"E73C",x"E73C",x"EF7E",x"E71C",x"AD54",x"62C8",x"3941",x"4120",
									 x"59C0",x"6241",x"7261",x"82A1",x"8AE1",x"9B21",x"A321",x"AB62",x"B382",x"BBA2",
									 x"BBC2",x"C3E2",x"C3E2",x"C3E2",x"C402",x"C402",x"C403",x"C402",x"C402",x"C423",
									 x"C403",x"BC02",x"BC02",x"BC02",x"B3E2",x"ABA2",x"AB82",x"9B42",x"9340",x"BCE4",
									 x"E6A6",x"F786",x"FFA6",x"FF66",x"FF26",x"FF05",x"FEE5",x"FEE5",x"FEC5",x"FEC5",
									 x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE45",x"FE24",x"FE05",
									 x"FDE4",x"FDC4",x"FD84",x"F543",x"F523",x"FCE3",x"F4A4",x"F4A6",x"E4CA",x"D551",
									 x"C5D6",x"BE17",x"C618",x"DEDB",x"EF3C",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",
									 x"FFBD",x"F6D8",x"F56D",x"EC66",x"EC02",x"F442",x"F483",x"F4C3",x"FCE3",x"FD04",
									 x"FD24",x"FD45",x"FD65",x"FD65",x"FDA5",x"FE08",x"FE6E",x"FF16",x"FF7A",x"FF7A",
									 x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FEEF",x"FEEF",x"FEEF",x"FECE",x"EE6C",x"BCC9",x"7282",x"5180",x"59A0",x"6A00",
									 x"7261",x"7A61",x"8281",x"8AA1",x"92E1",x"9B02",x"9B02",x"A322",x"A322",x"A342",
									 x"A342",x"AB42",x"AB42",x"AB42",x"AB42",x"AB42",x"AB42",x"A342",x"A342",x"A322",
									 x"A322",x"9B02",x"9B02",x"9B02",x"8AC1",x"7A40",x"7AC0",x"D629",x"FFCC",x"FFAB",
									 x"FF2A",x"FEA8",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE46",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE85",x"FEA5",x"FEC6",x"F665",x"D544",x"9B62",x"69A0",x"58E0",
									 x"5920",x"6160",x"6160",x"6160",x"69E2",x"938A",x"CDF5",x"DEBA",x"E71C",x"E71C",
									 x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"EF5D",
									 x"EF7E",x"E73C",x"C617",x"7B6B",x"3942",x"4100",x"51A0",x"6221",x"6A61",x"7AA1",
									 x"8AE1",x"9B01",x"9B21",x"AB62",x"B382",x"BBA2",x"BBC2",x"C3E2",x"C3E2",x"C3E2",
									 x"CC03",x"C402",x"C403",x"C403",x"C423",x"C422",x"C403",x"C403",x"C403",x"BC03",
									 x"BBE3",x"B3C2",x"ABA1",x"A362",x"9321",x"B464",x"CDA4",x"EF06",x"FFC7",x"FF86",
									 x"FF46",x"FF06",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",
									 x"FE85",x"FE85",x"FE65",x"FE45",x"FE24",x"FE04",x"FDE4",x"FDC4",x"FDA4",x"F543",
									 x"F543",x"FD03",x"F4A3",x"F485",x"ECA8",x"D52F",x"C5D5",x"BDF6",x"BDF8",x"D6BB",
									 x"E73C",x"F79D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FF7C",x"F675",x"ED0B",x"E425",
									 x"F402",x"F442",x"F483",x"F4C3",x"FCE4",x"FD04",x"FD44",x"FD64",x"FD64",x"FD84",
									 x"FDC6",x"FE4B",x"FEB1",x"FF37",x"FF7A",x"FF7A",x"FF79",x"FF79",x"FF79",x"FF78",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF35",
									 x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FEEF",x"FECE",
									 x"EE4C",x"BCC8",x"7282",x"5180",x"59A0",x"6A00",x"7261",x"7A61",x"8281",x"8AA1",
									 x"92E1",x"9302",x"9B02",x"A322",x"A322",x"A342",x"A342",x"AB42",x"AB42",x"AB42",
									 x"AB62",x"AB62",x"AB42",x"AB42",x"A342",x"A342",x"A322",x"9B22",x"9B22",x"9B22",
									 x"8AC1",x"7200",x"7A80",x"D629",x"FFCC",x"FFAB",x"FF2A",x"FEA8",x"FE67",x"FE67",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE66",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FEA5",
									 x"FEC5",x"FE86",x"DD85",x"A3A2",x"71C1",x"50E0",x"5900",x"6160",x"6180",x"6160",
									 x"6181",x"8B29",x"C5D5",x"DEDB",x"E71C",x"E71C",x"E73C",x"E73C",x"E73C",x"E73C",
									 x"E73C",x"E73C",x"EF5D",x"EF5D",x"E73C",x"EF5D",x"EF7D",x"EF5D",x"DEDA",x"942E",
									 x"3921",x"3900",x"51A0",x"6221",x"6A41",x"7A81",x"8AC1",x"9B01",x"9B21",x"AB62",
									 x"B382",x"BBA2",x"BBC2",x"C3E2",x"C3E2",x"C402",x"CC03",x"C403",x"C403",x"C403",
									 x"C423",x"C423",x"C423",x"C423",x"C423",x"BC03",x"BC02",x"B3E2",x"B3C2",x"AB82",
									 x"9B42",x"A3E2",x"AC62",x"DE44",x"FFA7",x"FFA6",x"FF66",x"FF26",x"FEE5",x"FEE5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",
									 x"FE24",x"FE04",x"FDE4",x"FDC4",x"FDA4",x"F563",x"F543",x"FD03",x"F4C3",x"F484",
									 x"EC87",x"D50D",x"CDB4",x"BDD6",x"BDD7",x"CE7A",x"DEFB",x"EF5D",x"FFDF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFDF",x"FF3A",x"F5F2",x"ECC9",x"EC24",x"F422",x"F462",x"F4A3",x"F4C3",
									 x"FCE4",x"FD04",x"FD44",x"FD64",x"FD84",x"F583",x"FDE7",x"FE8E",x"FEF4",x"FF58",
									 x"FF99",x"FF79",x"FF59",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FEEE",x"FECE",x"EE4C",x"C4E9",x"72A3",x"5180",
									 x"59A0",x"6A01",x"7241",x"7A61",x"8281",x"8AC1",x"92E1",x"9302",x"9B02",x"9B22",
									 x"A322",x"A342",x"A342",x"AB42",x"AB42",x"AB42",x"AB42",x"AB42",x"AB42",x"AB62",
									 x"A362",x"A342",x"A322",x"9B22",x"9B02",x"9302",x"8AC1",x"7A40",x"82E1",x"D629",
									 x"FFCC",x"FFAB",x"FF29",x"FEA7",x"FE67",x"FE47",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",x"FE86",x"FE86",x"FE65",
									 x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEA6",x"DDA4",x"ABE3",
									 x"7201",x"50C0",x"5900",x"6980",x"6180",x"6140",x"6161",x"8309",x"C5B5",x"D6DB",
									 x"E71C",x"E71C",x"E71C",x"E73C",x"E73C",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",
									 x"E73C",x"EF5D",x"EF7D",x"EF7D",x"EF5C",x"A4B1",x"3922",x"38E0",x"51A0",x"6221",
									 x"6A41",x"7A81",x"8AC1",x"9B02",x"9B22",x"AB62",x"B3A2",x"BBA2",x"BBC2",x"C3E2",
									 x"C3E2",x"C3E2",x"C403",x"C402",x"C422",x"C423",x"C422",x"C422",x"C423",x"C423",
									 x"C403",x"BC02",x"BC02",x"B402",x"B3C2",x"ABA3",x"A382",x"9B62",x"9BA1",x"CDC4",
									 x"FF67",x"FFA6",x"FF86",x"FF26",x"FF05",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",
									 x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE24",x"FE24",x"FE04",x"FDE4",
									 x"FDA4",x"F583",x"F543",x"FD03",x"FCC3",x"F4A3",x"EC85",x"DCEB",x"CD92",x"BDB5",
									 x"BDD7",x"CE59",x"D6BA",x"EF5C",x"FFBF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FEF8",x"F5B0",
									 x"EC88",x"EC24",x"F422",x"F462",x"F4A3",x"F4E3",x"FD04",x"FD24",x"FD44",x"FD64",
									 x"FD84",x"FD84",x"F609",x"FEB1",x"FF17",x"FF59",x"FF99",x"FF79",x"FF79",x"FF79",
									 x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FF11",
									 x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECF",
									 x"FEEE",x"FECE",x"F68C",x"CD29",x"82E4",x"5140",x"5140",x"6A01",x"7241",x"7A61",
									 x"82A2",x"8AC1",x"8AE1",x"92E2",x"9302",x"9B22",x"9B22",x"A342",x"A342",x"A342",
									 x"AB42",x"AB42",x"A342",x"A342",x"A342",x"A362",x"A342",x"A342",x"9B22",x"9B22",
									 x"9B02",x"92E2",x"8AA1",x"8AC1",x"9382",x"DE69",x"FFCC",x"FF8B",x"FF29",x"FEA7",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",
									 x"FE84",x"FEA5",x"FEA5",x"FEC6",x"E5E3",x"B443",x"7A22",x"50C0",x"58E0",x"6180",
									 x"61A0",x"6140",x"6141",x"82C9",x"C595",x"D6DB",x"E73C",x"E71C",x"E71C",x"E73C",
									 x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF7D",x"F77D",
									 x"F79E",x"AD13",x"3942",x"3100",x"49A0",x"6201",x"6A41",x"7281",x"82C1",x"9302",
									 x"9B22",x"AB62",x"B382",x"BBA2",x"BBC2",x"C3E2",x"C3E3",x"C3E3",x"C403",x"C403",
									 x"C422",x"C422",x"CC22",x"CC23",x"C422",x"C422",x"C403",x"C402",x"BC02",x"BC02",
									 x"B3C3",x"B3A2",x"AB82",x"9B42",x"9341",x"C524",x"F707",x"FFA6",x"FFC6",x"FF46",
									 x"FF05",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",
									 x"FE85",x"FE45",x"FE44",x"FE24",x"FE04",x"FDE4",x"FDC4",x"F583",x"F563",x"FD23",
									 x"FCE3",x"F4A2",x"EC84",x"DCC9",x"D570",x"BD94",x"BDB6",x"C639",x"D69A",x"E73C",
									 x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"FE96",x"F52D",x"EC66",x"EC03",x"F422",x"F463",
									 x"F4C3",x"F4E3",x"FD04",x"FD24",x"FD44",x"FD65",x"FD85",x"FDA5",x"F62B",x"FEF3",
									 x"FF39",x"FF7A",x"FF99",x"FF79",x"FF79",x"FF99",x"FF99",x"FF99",x"FF98",x"FF78",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF55",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FF11",x"FEF0",x"FEF0",x"FED0",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECF",x"FEEE",x"FEEE",x"FEAD",x"DDCC",
									 x"9BC7",x"5141",x"4940",x"61E1",x"7221",x"7A61",x"7A81",x"82A1",x"8AC1",x"92E2",
									 x"9302",x"9B02",x"9B22",x"9B22",x"A342",x"A342",x"A342",x"A342",x"A342",x"A342",
									 x"A342",x"A342",x"9B22",x"9B22",x"9B22",x"9B02",x"9302",x"8AA1",x"8281",x"9B63",
									 x"AC84",x"EF0A",x"FFCC",x"FF6B",x"FEE9",x"FE87",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FE84",x"FEA5",x"FEA5",x"FEE6",
									 x"E623",x"BC84",x"7A42",x"50C0",x"50E0",x"6160",x"61A0",x"6140",x"5921",x"82A8",
									 x"C595",x"D6FB",x"E73C",x"E71C",x"E71C",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",
									 x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF7D",x"F79D",x"FFDF",x"B575",x"41A4",x"3921",
									 x"4980",x"5A01",x"6241",x"7281",x"82C1",x"92E1",x"9B22",x"AB62",x"B382",x"BBA2",
									 x"BBC2",x"C3E2",x"C3E3",x"C3E3",x"C3E3",x"C403",x"C422",x"C422",x"CC22",x"CC22",
									 x"C422",x"C422",x"C423",x"C402",x"BC02",x"BC03",x"BBE4",x"B3C3",x"ABA2",x"9B21",
									 x"92E2",x"AC63",x"DE65",x"F785",x"FFC6",x"FF66",x"FF25",x"FEE5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE65",x"FE45",x"FE24",
									 x"FE24",x"FE04",x"FDE4",x"FDA4",x"FD83",x"FD24",x"FCE3",x"FCA2",x"F483",x"E4A8",
									 x"D50E",x"C593",x"BDB6",x"C5F8",x"CE79",x"DEFB",x"F77E",x"FFDF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF9C",
									 x"F634",x"F4CB",x"F445",x"EC03",x"F442",x"F483",x"F4C4",x"FCE4",x"FD04",x"FD24",
									 x"FD65",x"FD65",x"FD65",x"FDA7",x"FE4E",x"FF35",x"FF7A",x"FF7A",x"FF99",x"FF79",
									 x"FF79",x"FF99",x"FF99",x"FF99",x"FF98",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF55",x"FF55",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECF",x"FEEE",x"FEEE",x"FECD",x"F68D",x"B4A9",x"59A1",x"5140",x"59C1",
									 x"6A21",x"7241",x"7A61",x"82A2",x"8AC1",x"92C2",x"92E3",x"92E2",x"9B02",x"9B22",
									 x"9B22",x"A322",x"A322",x"A322",x"A322",x"A322",x"A342",x"9B22",x"9B22",x"9B22",
									 x"9B22",x"92E1",x"92C1",x"8260",x"7A81",x"AC45",x"CDC7",x"F76B",x"FFAB",x"FF4A",
									 x"FEC9",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE47",
									 x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",
									 x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEE6",x"EE64",x"BCA3",x"8262",x"48A0",
									 x"50E0",x"6160",x"61C0",x"6160",x"5920",x"7AA8",x"BD74",x"DEFB",x"E73C",x"E73C",
									 x"E73C",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",
									 x"EF7D",x"F79E",x"FFDF",x"BDB6",x"5206",x"4161",x"4980",x"59E0",x"6241",x"7261",
									 x"82C1",x"92E1",x"9B01",x"A342",x"B382",x"BBA2",x"BBC2",x"C3E3",x"C3E3",x"C3E2",
									 x"C403",x"C403",x"C422",x"C422",x"CC22",x"C422",x"C422",x"C422",x"C422",x"C422",
									 x"C422",x"BC03",x"BBE3",x"B3E3",x"B3C2",x"A342",x"9322",x"A3E2",x"CDA4",x"EF45",
									 x"FFC6",x"FFA6",x"FF46",x"FEE5",x"FEE5",x"FEE6",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE24",x"FE24",x"FE04",x"FDE4",x"FDA4",
									 x"FD84",x"FD44",x"FD03",x"F4C2",x"F483",x"E487",x"DCEC",x"C593",x"BDB6",x"BDF8",
									 x"C659",x"DEFB",x"F77D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF9B",x"FDF1",x"F489",x"F424",x"EC22",
									 x"F463",x"F4A3",x"F4C4",x"FD04",x"FD24",x"FD45",x"FD65",x"FD64",x"FD65",x"FDC9",
									 x"FE71",x"FF57",x"FF9A",x"FF7A",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",
									 x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FEEF",x"FEEE",
									 x"FECE",x"F6CD",x"C52A",x"7282",x"5980",x"5980",x"6201",x"7201",x"7A61",x"8282",
									 x"82A1",x"8AA2",x"8AC2",x"92E2",x"9B02",x"9B02",x"9B02",x"9B02",x"9B02",x"9B22",
									 x"9B22",x"9B22",x"9B21",x"9B21",x"9B02",x"9B22",x"9B01",x"92E1",x"92C2",x"8261",
									 x"82C1",x"B506",x"DE89",x"F76B",x"FF8A",x"FF09",x"FEA9",x"FE48",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE46",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FEA5",
									 x"FEA4",x"FF05",x"EE64",x"C4C3",x"8282",x"48A0",x"50C0",x"6160",x"61A0",x"5940",
									 x"5920",x"7AA8",x"BD74",x"DEDA",x"EF3D",x"E73C",x"E73C",x"EF5D",x"EF5C",x"EF5D",
									 x"EF7D",x"EF7D",x"EF7D",x"EF5D",x"EF5D",x"EF5D",x"EF7D",x"F79E",x"FFDF",x"C5D6",
									 x"5A67",x"4982",x"4980",x"59E0",x"6220",x"7241",x"82C2",x"8AE1",x"9B01",x"A342",
									 x"AB82",x"BBA2",x"BBC2",x"C3E3",x"C3E3",x"C3E2",x"C403",x"C403",x"C403",x"CC22",
									 x"CC22",x"C422",x"C422",x"C422",x"C422",x"C422",x"C423",x"BC22",x"BC02",x"B3E2",
									 x"B3E3",x"A362",x"9B42",x"9B82",x"BD04",x"EF07",x"FFC6",x"FFC6",x"FF67",x"FF05",
									 x"FEE6",x"FEC6",x"FEC6",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE65",
									 x"FE65",x"FE44",x"FE24",x"FE04",x"FDE4",x"FDA4",x"FD84",x"FD44",x"F503",x"F4C2",
									 x"F4A2",x"EC85",x"E4CA",x"D572",x"C5D6",x"BDF7",x"C639",x"DEDA",x"EF7D",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDF",x"FF5A",x"F56F",x"EC47",x"F403",x"F422",x"F463",x"F4A3",x"FCE4",x"FD04",
									 x"FD24",x"FD45",x"FD65",x"FD63",x"FD84",x"FDE9",x"FEB2",x"FF78",x"FF9A",x"FF7A",
									 x"FF79",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FEEE",x"FEEF",x"E60C",x"AC47",
									 x"8304",x"59A0",x"59A1",x"69E0",x"7220",x"7A61",x"82A1",x"82A1",x"8AC1",x"8AC1",
									 x"92E1",x"92E1",x"92E1",x"9B01",x"9B02",x"9B02",x"9B02",x"9B02",x"9B01",x"9B02",
									 x"9B02",x"9B02",x"92E2",x"8A81",x"7A20",x"7A60",x"9BC3",x"D629",x"F76C",x"FF8B",
									 x"FF29",x"FEE8",x"FE88",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",
									 x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA4",x"FF05",x"EE84",x"C504",
									 x"8AC2",x"50C0",x"50C0",x"6140",x"6980",x"6140",x"5100",x"7287",x"BD74",x"D6DA",
									 x"E73D",x"E73C",x"E73C",x"EF5D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",
									 x"EF7D",x"EF7D",x"EF7D",x"F79E",x"FFDF",x"CE17",x"6AE9",x"51E4",x"4160",x"51C0",
									 x"6220",x"7241",x"82A2",x"8AE1",x"9B01",x"A342",x"AB82",x"B3A2",x"BBC2",x"BBE3",
									 x"C3E3",x"C3E2",x"C403",x"C403",x"CC23",x"CC22",x"CC23",x"CC23",x"CC23",x"C423",
									 x"C423",x"C423",x"C423",x"BC23",x"BC02",x"BC02",x"B403",x"ABA2",x"A383",x"9321",
									 x"A442",x"DE66",x"F766",x"FFC6",x"FF86",x"FF26",x"FEE5",x"FEC5",x"FEC6",x"FEC5",
									 x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE65",x"FE45",x"FE24",x"FE24",
									 x"FDE4",x"FDA4",x"FD84",x"FD44",x"F523",x"F4E2",x"F4A2",x"EC85",x"E4A9",x"D551",
									 x"CDD5",x"B5D7",x"BE18",x"D69A",x"E73C",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFBD",x"FED8",x"ED2D",x"F446",
									 x"EC03",x"F443",x"F483",x"F4C3",x"FD04",x"FD25",x"FD45",x"FD45",x"FD65",x"FD83",
									 x"FD84",x"FE0A",x"FEF3",x"FF78",x"FF9A",x"FF9A",x"FF79",x"FF99",x"FF99",x"FF79",
									 x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FEEF",x"F6AE",x"E5EC",x"BCA8",x"7AA3",x"59A1",x"5980",
									 x"61A0",x"7221",x"7A61",x"8281",x"82A1",x"8AA1",x"8AC1",x"8AE1",x"92E1",x"92E1",
									 x"9301",x"9AE2",x"9AE2",x"92E1",x"92E1",x"92E2",x"92C2",x"92C2",x"8260",x"8240",
									 x"82A2",x"9BA4",x"CDA8",x"F72B",x"FFAB",x"FF6A",x"FEE8",x"FEA8",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE67",x"FE47",x"FE47",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE66",x"FE86",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FEA5",x"FEC4",x"FF05",x"F6C5",x"CD44",x"9303",x"5100",x"50C0",x"6140",
									 x"6980",x"6140",x"5100",x"7287",x"B554",x"D6DA",x"E73C",x"E71C",x"E73C",x"EF5D",
									 x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF9E",x"F77D",x"F79E",
									 x"FFDF",x"CE37",x"7B6B",x"5A25",x"4141",x"51A0",x"6220",x"6A40",x"82A2",x"8AE1",
									 x"9301",x"A342",x"AB82",x"B3A2",x"BBA2",x"BBE3",x"C3E2",x"C3E2",x"C403",x"C403",
									 x"CC23",x"CC23",x"CC23",x"CC23",x"CC23",x"C423",x"C422",x"C422",x"C423",x"C423",
									 x"BC22",x"BC02",x"B403",x"ABC2",x"ABA3",x"92E1",x"9BC2",x"CDC5",x"E6E5",x"FFC6",
									 x"FF86",x"FF46",x"FF05",x"FEC5",x"FEE6",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",
									 x"FEA5",x"FE85",x"FE85",x"FE45",x"FE24",x"FE25",x"FDE4",x"FDC4",x"FDA4",x"FD44",
									 x"FD24",x"F503",x"F4A3",x"EC84",x"E4A8",x"D52F",x"CD93",x"BDD6",x"BE18",x"CE79",
									 x"E71C",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFDE",x"FF7C",x"FE96",x"ECEB",x"F425",x"EC23",x"F463",x"F4A3",x"F4C3",
									 x"F4E4",x"FD24",x"FD24",x"FD45",x"FD85",x"FD84",x"F5A5",x"FE2B",x"FF15",x"FF79",
									 x"FF9A",x"FF7A",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FEEF",x"FECE",x"FECE",x"FEEF",
									 x"FEEE",x"F6AD",x"DDCA",x"A3C5",x"7241",x"61C0",x"61A0",x"69E1",x"7221",x"7A42",
									 x"7A62",x"8281",x"82A1",x"82A1",x"8AC1",x"8AC1",x"8AC2",x"8AC1",x"8AC1",x"8AC1",
									 x"92E1",x"8AC2",x"8AA2",x"8281",x"7A60",x"82C0",x"9B83",x"BCE6",x"E6A9",x"FF6A",
									 x"FF6A",x"FF09",x"FEC8",x"FE87",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE46",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE65",x"FE86",
									 x"FE85",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEC4",x"FF05",
									 x"F6C4",x"D584",x"9342",x"5920",x"50C0",x"6140",x"6960",x"6140",x"5120",x"6A66",
									 x"AD32",x"D6B9",x"E73C",x"E73C",x"E73C",x"EF5D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",
									 x"EF7D",x"EF7D",x"EF7D",x"F79E",x"F77E",x"F79E",x"FFDF",x"CE58",x"83CD",x"5A67",
									 x"4141",x"51A1",x"6200",x"6A40",x"82A2",x"8AE2",x"9301",x"A342",x"AB82",x"B382",
									 x"BBA2",x"BBC3",x"C3E2",x"C3E2",x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC23",
									 x"CC23",x"C423",x"C422",x"C422",x"C423",x"C423",x"BC22",x"BC22",x"BC03",x"B3E2",
									 x"ABC3",x"9B01",x"9B82",x"C525",x"DE65",x"FFC7",x"FFA6",x"FF86",x"FF25",x"FEE5",
									 x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE45",
									 x"FE24",x"FE25",x"FDE4",x"FDC4",x"FDA4",x"FD64",x"FD24",x"F503",x"F4C2",x"F484",
									 x"ECA7",x"DD2D",x"CD92",x"BDB5",x"C618",x"CE59",x"E71C",x"EF7D",x"FFDF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FF3B",x"FE54",
									 x"ECCA",x"F424",x"F423",x"F463",x"F4A3",x"F4C3",x"FD04",x"FD24",x"FD44",x"FD65",
									 x"FD85",x"FDA4",x"F5C6",x"FE4D",x"FF36",x"FF9A",x"FF9A",x"FF7A",x"FF99",x"FF9A",
									 x"FF99",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEED",x"F68C",x"DDAB",
									 x"AC06",x"8304",x"7241",x"59A0",x"5980",x"61C1",x"7201",x"7241",x"7A61",x"8281",
									 x"82A2",x"82A2",x"8AA2",x"82A1",x"82A1",x"8281",x"7A60",x"7220",x"7220",x"7A41",
									 x"82E1",x"AC24",x"CD87",x"E689",x"FF4A",x"FF49",x"FF09",x"FEC8",x"FE88",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE67",x"FE47",
									 x"FE47",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE65",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FEA5",x"FEC4",x"FF05",x"F6E5",x"D5A4",x"9B82",x"5940",
									 x"58E0",x"6141",x"6180",x"6160",x"5120",x"6A66",x"AD11",x"D699",x"E71C",x"E73D",
									 x"E73D",x"EF5D",x"EF7D",x"EF7D",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",
									 x"F79E",x"F79E",x"FFDF",x"D699",x"946F",x"6AA8",x"3921",x"49A1",x"5A00",x"6A40",
									 x"7AA1",x"8AC1",x"9301",x"A342",x"AB62",x"B382",x"BBA2",x"BBC3",x"C3E2",x"C3E2",
									 x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC23",x"CC23",x"C423",x"C423",x"C423",
									 x"C423",x"C423",x"C422",x"BC22",x"BC22",x"B3E2",x"B3C2",x"A321",x"A383",x"B484",
									 x"CDC4",x"FF87",x"FFA6",x"FF86",x"FF46",x"FF06",x"FEE5",x"FEE5",x"FEE5",x"FEC5",
									 x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE25",x"FDE4",x"FDC4",
									 x"FDA4",x"FD64",x"FD44",x"F503",x"FCC3",x"F483",x"EC86",x"E4EC",x"D571",x"BDB5",
									 x"BDF7",x"C658",x"DEDB",x"EF5D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FF19",x"FE12",x"EC88",x"EC03",x"EC22",x"F463",
									 x"F4A3",x"FCE3",x"FD04",x"FD44",x"FD45",x"FD65",x"FD85",x"FDA5",x"FDC8",x"FE8F",
									 x"FF58",x"FF9A",x"FF9A",x"FF7A",x"FF99",x"FF9A",x"FF99",x"FF79",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",
									 x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEED",x"FEED",x"FEAD",x"DDCA",x"C4E8",x"9BC5",x"7AA2",
									 x"6A21",x"7221",x"7201",x"7201",x"6A00",x"7220",x"7221",x"7221",x"7221",x"7A40",
									 x"7A40",x"7A60",x"7A80",x"7A81",x"82E2",x"9363",x"AC65",x"DE08",x"F6EA",x"FF2A",
									 x"FF4A",x"FF09",x"FEA8",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",
									 x"FE65",x"FE85",x"FE85",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",
									 x"FEC5",x"FF05",x"F6E5",x"DDC4",x"9BA2",x"6140",x"58E0",x"6120",x"6180",x"6160",
									 x"5120",x"6A45",x"ACD0",x"D698",x"E71C",x"EF5D",x"EF5D",x"EF5D",x"EF7D",x"F79D",
									 x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"FFDF",x"DEFA",
									 x"A4F2",x"732A",x"3921",x"49A1",x"5A00",x"6A40",x"7AA1",x"82C1",x"92E1",x"A342",
									 x"AB62",x"B382",x"BBA2",x"BBC2",x"C3E2",x"C403",x"C403",x"C403",x"CC23",x"CC23",
									 x"CC23",x"CC23",x"CC23",x"CC23",x"C423",x"C423",x"C423",x"C423",x"C422",x"BC22",
									 x"BC22",x"B402",x"B3C2",x"AB82",x"A363",x"A3C3",x"BD23",x"FF67",x"FFC6",x"FFA6",
									 x"FF46",x"FF06",x"FEE6",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",
									 x"FE85",x"FE65",x"FE45",x"FE25",x"FE04",x"FDC4",x"FDA4",x"FD84",x"FD44",x"FD23",
									 x"FCE3",x"F483",x"F485",x"E4CA",x"D54F",x"BD94",x"BDF7",x"C638",x"D6BA",x"EF5D",
									 x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBD",
									 x"F6D7",x"FDB0",x"F467",x"EC23",x"F422",x"FC83",x"F4A3",x"FCE4",x"FD04",x"FD44",
									 x"FD45",x"FD65",x"FD84",x"FDA6",x"FDEA",x"FE91",x"FF79",x"FF9A",x"FF9A",x"FF9A",
									 x"FF9A",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",
									 x"FF14",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FEAD",x"F68D",x"FECD",
									 x"FECD",x"FEEE",x"FECD",x"F6AD",x"DDCA",x"BCC7",x"A3E5",x"9365",x"82E3",x"7A82",
									 x"7221",x"6A00",x"61C0",x"61A0",x"69C0",x"7220",x"8281",x"8AE2",x"9363",x"A404",
									 x"B4C6",x"C567",x"E669",x"FF0A",x"FF2A",x"FF09",x"FEC8",x"FEA8",x"FE87",x"FE67",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE86",x"FE85",x"FE65",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEC5",x"FF05",x"FEC5",x"DDC3",
									 x"A3C2",x"6160",x"58E0",x"6140",x"6180",x"6160",x"5920",x"6A24",x"ACAF",x"D678",
									 x"E71C",x"EF5D",x"EF7D",x"EF7D",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",
									 x"F79E",x"F79E",x"F79E",x"F79E",x"FFDF",x"E71B",x"B554",x"7B6B",x"3101",x"49A1",
									 x"5A00",x"6A41",x"7A81",x"82C1",x"8B02",x"9B42",x"AB61",x"B382",x"B3A2",x"BBC2",
									 x"C3E2",x"C403",x"C403",x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"C443",x"C423",x"C423",x"BC23",x"BC23",x"BC03",x"B3E2",x"ABA2",
									 x"A362",x"9B42",x"B484",x"F748",x"FFC5",x"FFC6",x"FF65",x"FF26",x"FEE6",x"FEE5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE45",x"FE24",
									 x"FE05",x"FDE4",x"FDC4",x"FDA4",x"FD64",x"F523",x"FCE3",x"F4A3",x"F484",x"E4C9",
									 x"D52E",x"C594",x"BDF7",x"C618",x"D6BA",x"E73C",x"EF7D",x"FFDF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"F6B6",x"F56E",x"F446",x"F403",
									 x"F422",x"FC83",x"FCA3",x"FCE4",x"FD04",x"FD44",x"FD44",x"FD64",x"FD84",x"FDA6",
									 x"FE0B",x"FEB2",x"FF79",x"FF9A",x"FF9A",x"FF9A",x"FF9A",x"FF99",x"FF79",x"FF79",
									 x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",x"FF14",x"FF34",x"FF14",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FECD",x"FECD",x"FECD",x"FECD",
									 x"F68C",x"E5EA",x"CD49",x"BCC8",x"AC26",x"9BA4",x"9343",x"8B02",x"8B02",x"8AE2",
									 x"8B02",x"9322",x"9BA4",x"AC24",x"B4A5",x"CD45",x"DDE7",x"E648",x"F6EA",x"FF09",
									 x"FEE8",x"FEA8",x"FE88",x"FE67",x"FE67",x"FE47",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE47",x"FE47",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE86",x"FE85",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FEA5",x"FEA4",x"FF05",x"F6C5",x"E5E4",x"ABE2",x"6180",x"5900",x"6140",
									 x"6180",x"6160",x"5920",x"6A24",x"A46E",x"CE37",x"DEFB",x"EF5D",x"EF7D",x"EF7D",
									 x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",
									 x"FFDF",x"EF3C",x"C5D6",x"83AD",x"3102",x"49A1",x"5A01",x"6A41",x"7A81",x"82C1",
									 x"8B02",x"9B42",x"AB61",x"B382",x"B3A2",x"BBC2",x"C3E2",x"C403",x"C403",x"C403",
									 x"C403",x"CC23",x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C423",
									 x"C423",x"C423",x"BC23",x"B402",x"B3E2",x"B3C2",x"A362",x"9301",x"AC43",x"EF07",
									 x"FFC6",x"FFC6",x"FF66",x"FF26",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE45",x"FE24",x"FE05",x"FDE4",x"FDC4",x"FDA4",
									 x"FD64",x"FD23",x"FD03",x"F4C3",x"F484",x"ECA8",x"D50D",x"C593",x"BDD6",x"C617",
									 x"CE99",x"E71C",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFE",x"F77B",x"F654",x"F50C",x"F425",x"F402",x"F442",x"FC83",x"FCC4",x"FCE4",
									 x"FD04",x"FD44",x"FD44",x"FD64",x"FD84",x"FDC7",x"FE2C",x"FEF4",x"FF79",x"FF9A",
									 x"FF7A",x"FF9A",x"FF9A",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",
									 x"FF34",x"FF34",x"FF14",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEEC",x"FEED",x"FEED",x"FEAC",x"F66C",
									 x"EE2A",x"DDC9",x"D588",x"D567",x"D546",x"D546",x"D546",x"D587",x"DDC7",x"E608",
									 x"EE89",x"FEC9",x"FF09",x"FF09",x"FF09",x"FEA8",x"FE87",x"FE67",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE86",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA4",x"FF05",
									 x"F6C4",x"E624",x"B443",x"69C0",x"5920",x"5940",x"6180",x"6140",x"5920",x"6A23",
									 x"9C2D",x"CE16",x"DEDB",x"EF5D",x"EF7D",x"F79E",x"F79E",x"F79E",x"F7BE",x"F7BE",
									 x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"FFDF",x"F77D",x"D638",x"8BEF",
									 x"3902",x"4161",x"5A01",x"6A41",x"7281",x"82C1",x"8AE2",x"9B22",x"AB61",x"B382",
									 x"B3A2",x"BBC2",x"C3C2",x"C3E3",x"C403",x"C403",x"C403",x"CC23",x"CC23",x"CC23",
									 x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",x"C442",x"C443",x"C443",x"BC23",x"BC03",
									 x"B402",x"B3E2",x"A362",x"9301",x"A402",x"E686",x"F786",x"FFC6",x"FF66",x"FF46",
									 x"FF05",x"FEE5",x"FEC5",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE65",
									 x"FE65",x"FE45",x"FE25",x"FDE4",x"FDC4",x"FDA4",x"FD64",x"FD23",x"FD03",x"F4C3",
									 x"F484",x"ECA7",x"D4EC",x"CD72",x"C5D5",x"BDF7",x"CE79",x"DEFB",x"EF7D",x"F7BE",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"F719",x"F5F2",x"F4CA",
									 x"F425",x"F422",x"F463",x"F4A3",x"FCC4",x"FD04",x"FD24",x"FD44",x"FD64",x"FD84",
									 x"FD85",x"FDE8",x"FE6E",x"FEF5",x"FF9A",x"FF9A",x"FF7A",x"FF7A",x"FF7A",x"FF99",
									 x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",x"FF14",x"FF34",
									 x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",
									 x"FEF1",x"FF11",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FECD",x"FECD",
									 x"FEAD",x"FEAC",x"FEAB",x"FECC",x"FECC",x"FECB",x"FECB",x"FEAA",x"F689",x"F688",
									 x"FE88",x"FE88",x"FE88",x"F6A7",x"F6C7",x"FEC8",x"FEA8",x"FEA8",x"FEA8",x"FEA8",
									 x"FE87",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",
									 x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE47",
									 x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA4",x"FF05",x"FEC5",x"EE44",x"BC83",x"7200",
									 x"5940",x"5920",x"6160",x"6160",x"5940",x"6A02",x"9C0B",x"CDD5",x"DEDB",x"EF5D",
									 x"EF7D",x"F79E",x"F79E",x"F79E",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",
									 x"F7BE",x"F7BE",x"FFDF",x"F79E",x"DEBA",x"9450",x"3102",x"4161",x"59E0",x"6221",
									 x"7281",x"82C1",x"8AE2",x"9B22",x"AB41",x"B382",x"B3A2",x"BBC2",x"C3C2",x"C3E3",
									 x"C403",x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",
									 x"CC43",x"C442",x"C442",x"C443",x"BC43",x"BC23",x"B402",x"B3E2",x"A362",x"9B01",
									 x"A3C2",x"D5E5",x"F746",x"FFC7",x"FF86",x"FF46",x"FF05",x"FEE5",x"FEC5",x"FEE5",
									 x"FEE5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE45",x"FE25",x"FE05",
									 x"FDE4",x"FDC4",x"FD84",x"F543",x"FD23",x"F4C3",x"F483",x"EC86",x"DCEB",x"CD71",
									 x"C5B4",x"BDD6",x"CE79",x"DEFB",x"EF5D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFBD",x"F6D7",x"F5B0",x"F4A9",x"F424",x"F422",x"F463",x"F4A3",
									 x"FCE4",x"FD04",x"FD24",x"FD44",x"FD64",x"FD85",x"F585",x"FDE8",x"FE6E",x"FF16",
									 x"FF9A",x"FF9A",x"FF7A",x"FF7A",x"FF7A",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",
									 x"FF55",x"FF34",x"FF34",x"FF34",x"FF14",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FF11",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FECC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FECC",x"FECB",x"FECA",x"FEC9",x"FEC8",x"FEC8",x"FEC8",x"FEE8",
									 x"FEE7",x"FEC8",x"FE87",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",
									 x"FEA4",x"FF05",x"FEC5",x"EE64",x"BCA3",x"7A41",x"6140",x"5920",x"5960",x"6160",
									 x"5940",x"61E1",x"93CA",x"CDD4",x"DEDA",x"EF5D",x"EF7D",x"F79E",x"F79E",x"F7BE",
									 x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"FF9E",x"FFBF",x"FFDF",x"FFDF",
									 x"EF1B",x"9C71",x"3102",x"4140",x"51E0",x"6220",x"7281",x"82A1",x"8AE1",x"9B22",
									 x"AB41",x"B362",x"B3A2",x"BBC2",x"C3C2",x"C3E3",x"C403",x"C403",x"C403",x"CC23",
									 x"CC23",x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",x"C442",x"C442",x"C443",
									 x"BC43",x"BC23",x"B422",x"B3E2",x"AB82",x"9B22",x"A3A2",x"CD64",x"EF06",x"FFC7",
									 x"FFA6",x"FF66",x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEA5",x"FEA5",
									 x"FEA5",x"FE85",x"FE65",x"FE45",x"FE25",x"FE05",x"FDE4",x"FDC4",x"FD83",x"FD43",
									 x"FD23",x"F4C3",x"F4A3",x"F485",x"DCCA",x"CD50",x"C593",x"BDB5",x"C659",x"DEDB",
									 x"E73C",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF9D",x"F676",
									 x"F56E",x"F488",x"F424",x"F443",x"F463",x"F4A3",x"FCE4",x"FD04",x"FD24",x"FD64",
									 x"FD65",x"FD85",x"F585",x"FDE8",x"FE8F",x"FF36",x"FF7A",x"FF9A",x"FF7A",x"FF7A",
									 x"FF79",x"FF99",x"FF99",x"FF79",x"FF79",x"FF99",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FEF2",x"FEF1",x"FEF1",x"FF11",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAC",x"FEAD",x"FECC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8B",
									 x"FE6A",x"FE68",x"FE67",x"FE67",x"FE88",x"FE88",x"FE87",x"FE67",x"FE67",x"FE46",
									 x"FE46",x"FE47",x"FE47",x"FE67",x"FE68",x"FE48",x"FE68",x"FE67",x"FE47",x"FE47",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA4",x"FF05",x"FEC5",x"EE64",
									 x"C4C3",x"7A40",x"6140",x"5920",x"5940",x"6160",x"6140",x"61C0",x"93A9",x"CDD4",
									 x"DEBA",x"EF5D",x"EF7D",x"F79E",x"F79E",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",
									 x"F7BE",x"F7BE",x"F79E",x"F7BF",x"FFDF",x"FFDF",x"F75C",x"A4B1",x"3922",x"4140",
									 x"51E0",x"6200",x"7261",x"7AA1",x"8AC1",x"9B22",x"AB41",x"AB82",x"B3A2",x"BBC2",
									 x"C3E2",x"C3E3",x"C403",x"C403",x"C403",x"CC23",x"CC23",x"C423",x"CC23",x"CC43",
									 x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C443",x"C443",x"BC22",x"BC22",x"B402",
									 x"AB82",x"A342",x"A3A2",x"BCE3",x"E6C6",x"FFC7",x"FFA6",x"FF66",x"FF25",x"FEE5",
									 x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE45",
									 x"FE25",x"FE05",x"FDE4",x"FDC4",x"FD84",x"FD43",x"FD23",x"F4E3",x"F4A3",x"F485",
									 x"E4C9",x"D52E",x"C573",x"BD95",x"C639",x"D6BA",x"E71C",x"F79E",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F79C",x"F613",x"F50C",x"EC68",x"F403",x"F443",
									 x"F482",x"F4C3",x"FCE4",x"FD04",x"FD24",x"FD65",x"FD85",x"FD84",x"FD64",x"FE0A",
									 x"FED1",x"FF57",x"FF79",x"FF7A",x"FF7A",x"FF7A",x"FF79",x"FF99",x"FF79",x"FF79",
									 x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FE8B",x"FE8B",x"FE6A",x"FE49",x"FE47",x"FE46",x"FE46",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FEA5",x"FEA5",x"FEE5",x"FEE5",x"F684",x"C4E3",x"7A40",x"6140",x"5920",
									 x"5940",x"6160",x"6140",x"69A0",x"9369",x"C5B3",x"DEBA",x"EF5D",x"EF7D",x"EF7D",
									 x"F7BE",x"F7BF",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"FFBE",x"FFBE",
									 x"F7DF",x"FFDE",x"F79D",x"A512",x"3942",x"4140",x"51C0",x"6200",x"7262",x"82C2",
									 x"8AC2",x"9B22",x"A362",x"AB62",x"B3A2",x"BBC2",x"C3E2",x"C3E3",x"C403",x"C403",
									 x"C403",x"CC23",x"C423",x"C423",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",
									 x"C443",x"C443",x"C423",x"BC22",x"BC02",x"B403",x"ABA3",x"A381",x"9B82",x"AC63",
									 x"DE65",x"FFA7",x"FFC6",x"FF85",x"FF26",x"FEE6",x"FEE5",x"FEE5",x"FEE5",x"FEC5",
									 x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE45",x"FE45",x"FE05",x"FDE4",x"FDC4",
									 x"FDA4",x"FD43",x"FD24",x"F4E4",x"F4A4",x"ECA5",x"E4C7",x"DD2C",x"C572",x"B595",
									 x"C618",x"D6BA",x"E71C",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"F77C",x"F5F2",x"ECEC",x"EC47",x"F423",x"F443",x"F483",x"FCC3",x"FCE4",x"FD04",
									 x"FD24",x"FD64",x"FD65",x"FD64",x"FD85",x"FE2A",x"FEF2",x"FF58",x"FF79",x"FF7A",
									 x"FF79",x"FF9A",x"FF99",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",
									 x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8B",
									 x"FE8B",x"FE8A",x"FE69",x"FE47",x"FE46",x"FE47",x"FE67",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEE5",
									 x"FEE5",x"F685",x"CCE3",x"8260",x"6160",x"5920",x"6140",x"6160",x"6140",x"61A0",
									 x"8B68",x"C5B3",x"D6BA",x"EF5D",x"F79D",x"F79E",x"F79E",x"F7BF",x"F7BE",x"F7BE",
									 x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"FFDE",x"FFBE",x"FFDF",x"FFFF",x"F7BE",x"AD33",
									 x"4163",x"4140",x"51A0",x"6200",x"7261",x"7AC1",x"8AC2",x"9302",x"A341",x"AB62",
									 x"B382",x"BBC2",x"C3E2",x"C3E3",x"C403",x"C403",x"C403",x"CC23",x"C423",x"C423",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C443",x"C423",x"BC22",
									 x"BC22",x"B403",x"B3C3",x"A3A1",x"9B62",x"A402",x"DE45",x"FF87",x"FFA6",x"FF86",
									 x"FF46",x"FF06",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",
									 x"FE85",x"FE65",x"FE45",x"FE05",x"FDE4",x"FDC4",x"FDA4",x"FD63",x"FD24",x"F4E4",
									 x"F4C4",x"ECA5",x"ECC7",x"DD0C",x"C551",x"B595",x"BE18",x"CE79",x"DEFB",x"EF7D",
									 x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF7C",x"F5B0",x"F4EB",x"EC46",
									 x"F423",x"F463",x"F4A3",x"F4C3",x"FCE4",x"FD04",x"FD24",x"FD44",x"FD65",x"FD64",
									 x"FD85",x"FE2B",x"FF14",x"FF79",x"FF7A",x"FF7A",x"FF79",x"FF99",x"FF99",x"FF99",
									 x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8A",x"FE69",x"FE47",
									 x"FE47",x"FE47",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEC5",x"FEE5",x"F685",x"CD03",x"8260",
									 x"6160",x"5900",x"6140",x"6160",x"6160",x"69A0",x"8B68",x"C5B3",x"D6BA",x"EF7D",
									 x"F79E",x"F79E",x"F79E",x"F7BF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",
									 x"FFDF",x"FFBF",x"FFDF",x"FFFF",x"F7BE",x"AD54",x"41A3",x"3940",x"49A0",x"5A00",
									 x"7261",x"7AA1",x"82C2",x"9302",x"A341",x"AB62",x"B382",x"BBC2",x"BBE2",x"C3E2",
									 x"C403",x"C403",x"C403",x"CC23",x"CC23",x"C423",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"CC43",x"C443",x"C443",x"C443",x"C423",x"BC22",x"BC22",x"B403",x"B3C3",x"A3A2",
									 x"9B62",x"9BC2",x"DE25",x"F767",x"FFA6",x"FFA6",x"FF46",x"FF06",x"FEE5",x"FEE5",
									 x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE05",
									 x"FE04",x"FDC4",x"FDA4",x"FD84",x"FD44",x"F504",x"F4C3",x"ECA5",x"ECA6",x"E4EB",
									 x"CD30",x"BD95",x"BDF7",x"CE59",x"DEDB",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FF5B",x"F58F",x"F4C9",x"EC45",x"F422",x"F463",x"F483",x"FCC3",
									 x"FCE4",x"FD04",x"FD44",x"FD64",x"FD65",x"FD64",x"FDA6",x"FE4D",x"FF15",x"FF7A",
									 x"FF9A",x"FF79",x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",
									 x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",
									 x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FEF0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",
									 x"FEAC",x"FE8C",x"FE8B",x"FE6A",x"FE68",x"FE47",x"FE46",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",
									 x"FEC5",x"FEC5",x"FEE5",x"F6A5",x"CD03",x"8280",x"6160",x"5900",x"6140",x"6160",
									 x"6160",x"69A0",x"8B68",x"BDB3",x"D6BA",x"EF7D",x"F79E",x"F79E",x"F7BE",x"F7BF",
									 x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFBF",x"FFFF",x"FFFF",
									 x"F7BE",x"B554",x"49C4",x"3940",x"49A0",x"5A00",x"6A61",x"7AA1",x"82C2",x"9302",
									 x"A341",x"AB62",x"B382",x"BBC2",x"BBE2",x"C3E2",x"C403",x"CC03",x"C403",x"CC23",
									 x"CC23",x"C423",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C443",
									 x"C423",x"BC22",x"BC22",x"BC23",x"B3E3",x"ABA2",x"9B42",x"9BA1",x"D5C5",x"F767",
									 x"FFC7",x"FFA6",x"FF46",x"FF26",x"FF05",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE25",x"FE05",x"FDC4",x"FDA4",x"FD83",
									 x"FD43",x"F503",x"F4C3",x"F4A4",x"EC86",x"E4CA",x"CD0F",x"BD94",x"BDF7",x"CE59",
									 x"DEDB",x"EF5D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF3A",x"F54E",
									 x"EC88",x"EC24",x"FC22",x"F463",x"F4A3",x"FCC3",x"FD04",x"FD04",x"FD44",x"FD65",
									 x"FD85",x"FD85",x"FDC7",x"FE6E",x"FF36",x"FF7A",x"FF9A",x"FF79",x"FF99",x"FF99",
									 x"FF99",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",
									 x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FF12",x"FEF1",x"FEF1",x"FF11",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FEF0",x"FECF",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FE8C",x"FE8B",x"FE69",
									 x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEC5",x"FEC5",x"FEE6",x"FEA5",
									 x"D523",x"8280",x"6160",x"5900",x"6140",x"6160",x"6160",x"69A0",x"8B48",x"BDB3",
									 x"D6BA",x"EF7D",x"F79E",x"F79E",x"F7BF",x"F7DF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFBE",x"B574",x"49C4",x"4160",
									 x"49A0",x"5A00",x"6A61",x"7AA1",x"82C2",x"9302",x"A341",x"AB62",x"B382",x"BBC2",
									 x"BBE2",x"C3E2",x"C403",x"CC03",x"C403",x"CC23",x"CC23",x"C423",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"C443",x"C443",x"C443",x"C443",x"C443",x"BC23",x"BC42",x"BC23",
									 x"B3E3",x"ABC2",x"9B42",x"9B61",x"CD84",x"EF27",x"FFC7",x"FFA6",x"FF46",x"FF26",
									 x"FF05",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",
									 x"FE45",x"FE25",x"FE05",x"FDC5",x"FDA4",x"F584",x"F563",x"F503",x"F4C3",x"F484",
									 x"EC85",x"E4C9",x"CD0F",x"BD94",x"BDF7",x"C638",x"D6BA",x"EF5D",x"F7BE",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFE",x"FFFF",x"FF1A",x"F52D",x"EC67",x"EC04",x"FC22",x"F463",
									 x"F4A3",x"FCE4",x"FD04",x"FD04",x"FD44",x"FD64",x"FD65",x"FD85",x"FDE8",x"FE8F",
									 x"FF36",x"FF7B",x"FF9A",x"FF79",x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",
									 x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FE8C",x"FEAC",x"FE8C",x"FE8B",x"FE69",x"FE68",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FEA5",x"FEA5",x"FEC5",x"FEE5",x"FEC5",x"D544",x"82A1",x"6161",x"5100",
									 x"6140",x"6160",x"6160",x"61A0",x"8B48",x"BD93",x"D6BA",x"EF7D",x"F79E",x"F79E",
									 x"F7BF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",
									 x"FFFF",x"FFFF",x"FFBE",x"B574",x"49E4",x"4161",x"49A0",x"5A00",x"6A61",x"7AA1",
									 x"82C2",x"9302",x"A341",x"AB62",x"B382",x"BBC2",x"BBE2",x"C3E2",x"C403",x"C403",
									 x"C403",x"CC23",x"CC23",x"C423",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",
									 x"C443",x"C443",x"C443",x"C443",x"BC43",x"BC23",x"B3E3",x"ABC2",x"9B42",x"9341",
									 x"CD64",x"EF06",x"FFA7",x"FFA6",x"FF66",x"FF26",x"FF05",x"FEE5",x"FEE5",x"FEC5",
									 x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE25",x"FE05",x"FDC5",
									 x"FDC4",x"F5A4",x"F563",x"F523",x"F4C3",x"F483",x"EC84",x"E4A8",x"CD0E",x"BD74",
									 x"BDD7",x"C638",x"D6BA",x"E73C",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FF19",x"F50C",x"F446",x"EC04",x"F402",x"F463",x"F4A3",x"FCE4",x"FD04",x"FD04",
									 x"FD44",x"FD64",x"FD64",x"FDA5",x"FE09",x"FE90",x"FF37",x"FF7A",x"FF9A",x"FF7A",
									 x"FF99",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",
									 x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FED0",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FEAC",
									 x"FE8B",x"FE69",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEC5",
									 x"FEC5",x"FEC5",x"D544",x"82C1",x"6161",x"5100",x"6140",x"6160",x"6160",x"69A0",
									 x"8B28",x"C593",x"D6BA",x"F79D",x"F7BE",x"F7BE",x"F7BE",x"FFFF",x"FFDF",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"BD95",
									 x"5205",x"4161",x"49A0",x"5A00",x"7261",x"7AA1",x"82C2",x"9322",x"A361",x"AB82",
									 x"B382",x"BBC2",x"C3C2",x"C3E2",x"C403",x"C403",x"C402",x"CC22",x"CC22",x"CC23",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C443",x"C443",x"C443",
									 x"BC23",x"BC23",x"BBE2",x"B3C3",x"A362",x"9B41",x"CD25",x"E6A6",x"FF87",x"FFA6",
									 x"FF66",x"FF26",x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FE85",x"FE65",x"FE45",x"FE24",x"FE04",x"FDC5",x"FDC4",x"FD84",x"FD63",x"FD03",
									 x"F4C3",x"F4A3",x"F483",x"E4A7",x"CD0D",x"BD93",x"BDD7",x"C638",x"D69A",x"E73C",
									 x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FEF9",x"ECEB",x"F425",x"EBE3",
									 x"F402",x"FC83",x"F4A3",x"FCE4",x"FD04",x"FD24",x"FD44",x"FD64",x"FD64",x"FD85",
									 x"FE09",x"FE90",x"FF37",x"FF7A",x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",
									 x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FEAC",x"FE8B",x"FE69",x"FE48",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEC5",x"FEC5",x"FEC5",x"D564",x"8AE1",
									 x"6161",x"50E0",x"6140",x"6160",x"6160",x"69A0",x"8B27",x"C593",x"DEBA",x"F79D",
									 x"F7BE",x"F7BE",x"F7DF",x"FFFF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"BDB5",x"5245",x"3961",x"4180",x"5A00",
									 x"6A61",x"7A81",x"82C1",x"9302",x"9B41",x"AB62",x"B382",x"BBA2",x"C3C2",x"C3E2",
									 x"C403",x"C403",x"CC22",x"CC22",x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C443",x"C443",x"BC23",x"BC02",x"B3C3",
									 x"A362",x"9B41",x"C504",x"DE65",x"FF67",x"FFC6",x"FF86",x"FF46",x"FF05",x"FEE5",
									 x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE45",x"FE24",
									 x"FE04",x"FDE5",x"FDC4",x"FDA4",x"FD64",x"FD23",x"F4C3",x"F4A3",x"F483",x"E4A6",
									 x"D50D",x"BD94",x"BDD7",x"C618",x"D69A",x"E71C",x"F79E",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FEF8",x"ECAA",x"F405",x"EBE3",x"F422",x"F483",x"F4C3",x"F4E4",
									 x"FD04",x"FD24",x"FD44",x"FD64",x"FD64",x"FD85",x"FE2A",x"FEB1",x"FF37",x"FF9A",
									 x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF79",
									 x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",
									 x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECE",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",
									 x"FEAC",x"FEAC",x"FE8B",x"FE69",x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FEA4",x"FEC5",x"FEC5",x"FEC5",x"DD84",x"8AE1",x"6181",x"50E0",x"5940",x"6180",
									 x"6160",x"6180",x"8B07",x"C593",x"D6BA",x"F79D",x"F7BE",x"F7BE",x"F7DF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFBE",x"BDB6",x"5A66",x"4181",x"4180",x"59E0",x"6A61",x"7281",x"82C2",x"9302",
									 x"9B41",x"AB62",x"B382",x"BBC2",x"C3C2",x"C3E2",x"C403",x"CC03",x"CC22",x"CC22",
									 x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"C443",x"C443",x"C443",x"BC23",x"BC02",x"B3C3",x"A382",x"9B61",x"BCC3",x"D625",
									 x"F767",x"FFC7",x"FF86",x"FF46",x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE45",x"FE24",x"FE04",x"FDE5",x"FDC4",x"FDA4",
									 x"FD64",x"FD23",x"FCC3",x"F4A3",x"F463",x"E486",x"D50D",x"C593",x"BDD7",x"BDF8",
									 x"CE79",x"E71C",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FEF8",x"ECA9",
									 x"F404",x"EC03",x"FC22",x"F483",x"F4C3",x"F4E4",x"FD04",x"FD24",x"FD64",x"FD64",
									 x"FD64",x"FD85",x"FE0A",x"FEB1",x"FF37",x"FF9A",x"FF9A",x"FF9A",x"FF99",x"FF99",
									 x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",
									 x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FEAC",x"FE8B",x"FE69",
									 x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEC5",x"FEC5",x"FEE5",
									 x"DDA4",x"9301",x"69A1",x"50E0",x"6140",x"6181",x"6160",x"6180",x"8307",x"C572",
									 x"D6BA",x"F79D",x"F7BE",x"F7BE",x"F7DF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"C5D6",x"6287",x"4181",
									 x"4180",x"59E0",x"6A61",x"7281",x"82A2",x"9302",x"9B41",x"A362",x"B382",x"BBC2",
									 x"C3E2",x"C3E2",x"C403",x"C403",x"CC22",x"CC22",x"CC23",x"CC23",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C443",x"BC23",
									 x"BBE2",x"B3C3",x"A383",x"9B61",x"BCA3",x"D604",x"F767",x"FFC7",x"FF86",x"FF46",
									 x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FE85",
									 x"FE45",x"FE24",x"FE04",x"FDE5",x"FDC4",x"FDA4",x"FD64",x"FD23",x"FCC3",x"F4A3",
									 x"F463",x"EC86",x"D4EC",x"C593",x"BDD7",x"BE18",x"D699",x"E71C",x"F79E",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FED7",x"EC88",x"F404",x"EC03",x"FC22",x"F483",
									 x"F4C3",x"F4E4",x"FD04",x"FD24",x"FD64",x"FD64",x"FD64",x"FD86",x"FE2B",x"FED2",
									 x"FF58",x"FF9A",x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",
									 x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FE8C",x"FEAC",x"FEAC",x"FE8B",x"FE69",x"FE68",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FEA5",x"FEC5",x"FEE5",x"FEE5",x"DDA4",x"9301",x"69A1",x"50E0",
									 x"5940",x"6181",x"6160",x"6160",x"82E6",x"BD72",x"D6B9",x"F79D",x"F7BE",x"F7BE",
									 x"F7DF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFBE",x"C5F6",x"62C8",x"4182",x"4160",x"59E1",x"6A61",x"7281",
									 x"82A2",x"9301",x"9B41",x"A362",x"B382",x"BBC2",x"C3E2",x"C3E2",x"C403",x"C403",
									 x"CC22",x"CC22",x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"C443",x"C443",x"C443",x"BC23",x"BC02",x"B3C3",x"A383",x"9B61",
									 x"B483",x"CDE4",x"F747",x"FFA7",x"FF87",x"FF46",x"FF05",x"FEE5",x"FEE5",x"FEE5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE45",x"FE24",x"FE04",x"FDE5",
									 x"FDC4",x"FDA4",x"FD64",x"FD23",x"FCC3",x"F4A3",x"F463",x"EC65",x"D4EC",x"C573",
									 x"BDD7",x"BDF8",x"CE79",x"E71C",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FED7",x"EC68",x"F403",x"EBE3",x"F422",x"F483",x"F4C3",x"F4E4",x"FD04",x"FD24",
									 x"FD64",x"FD64",x"FD64",x"FD86",x"FE2B",x"FED2",x"FF58",x"FFBA",x"FF9A",x"FF9A",
									 x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FEAC",
									 x"FE8B",x"FE89",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEC5",
									 x"FEC5",x"FF05",x"DDC4",x"9321",x"69A1",x"50E0",x"5940",x"6181",x"6160",x"6160",
									 x"82C6",x"BD52",x"D6B9",x"F79D",x"F7BE",x"F7BE",x"F7DF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"C5F7",
									 x"6AC8",x"4182",x"4160",x"59E1",x"6A61",x"7A81",x"82A1",x"9301",x"9B41",x"A362",
									 x"B382",x"BBC2",x"C3C2",x"C3E2",x"C403",x"C403",x"CC22",x"CC22",x"CC23",x"CC23",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",
									 x"C443",x"BC23",x"BC02",x"B3E3",x"AB83",x"9B61",x"B483",x"CDC4",x"F747",x"FFC7",
									 x"FF87",x"FF46",x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FE85",x"FE85",x"FE45",x"FE24",x"FE04",x"FDE5",x"FDC4",x"FDA4",x"FD64",x"FD23",
									 x"F4C3",x"F4A3",x"F462",x"EC65",x"D4EB",x"C573",x"BDD7",x"BDF7",x"CE79",x"DEFB",
									 x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FED7",x"F447",x"F402",x"F3E2",
									 x"F442",x"F483",x"F4C3",x"F4E4",x"FD04",x"FD24",x"FD44",x"FD64",x"FD64",x"FD86",
									 x"FE2C",x"FED3",x"FF58",x"FF9A",x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",
									 x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAB",x"FE8B",x"FE89",x"FE68",x"FE47",
									 x"FE47",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEA5",x"FEC5",x"FEC5",x"FF05",x"DDC4",x"9321",
									 x"69A1",x"50E0",x"5940",x"6180",x"6180",x"6140",x"82A7",x"BD32",x"D699",x"F79D",
									 x"F7BE",x"F7DE",x"F7DF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"C617",x"6AC8",x"4182",x"4160",x"59E0",
									 x"6A61",x"7A81",x"82A1",x"9301",x"9B41",x"A362",x"B382",x"BBC2",x"C3C3",x"C3E3",
									 x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C443",x"BC23",x"BC02",x"B3E3",
									 x"AB83",x"9B61",x"B483",x"CDC4",x"F747",x"FFC7",x"FF86",x"FF46",x"FF05",x"FEE5",
									 x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE24",
									 x"FE04",x"FE05",x"FDC4",x"FDA4",x"FD64",x"FD23",x"F4E3",x"F4A3",x"F462",x"EC64",
									 x"D4CB",x"C573",x"B5D7",x"BDF7",x"CE79",x"E71C",x"F79E",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FED7",x"F447",x"EBE2",x"F3E2",x"F442",x"F483",x"F4C3",x"F4E4",
									 x"FD04",x"FD24",x"FD44",x"FD64",x"FD64",x"FD86",x"FE2C",x"FED3",x"FF58",x"FF7A",
									 x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",
									 x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAB",x"FE8A",x"FE89",x"FE68",x"FE47",x"FE47",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",
									 x"FEA5",x"FEC5",x"FEE5",x"FF05",x"E5C4",x"9321",x"69A1",x"50E0",x"5940",x"6180",
									 x"6180",x"6140",x"7A86",x"BD32",x"D6B9",x"F79D",x"F7DE",x"F7DE",x"F7DF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFBE",x"CE17",x"6AE9",x"4182",x"4160",x"59C0",x"6A41",x"7A61",x"82A1",x"9301",
									 x"9B41",x"A362",x"B382",x"BBA2",x"C3C3",x"C3E3",x"C403",x"C403",x"CC23",x"CC23",
									 x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"C443",x"C443",x"C423",x"BC23",x"BC02",x"B3E3",x"ABA3",x"9B61",x"B483",x"CDA4",
									 x"EF26",x"FFC7",x"FF86",x"FF46",x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE24",x"FE04",x"FE05",x"FDC4",x"FDA4",
									 x"FD84",x"FD24",x"F4E3",x"F4A3",x"F462",x"EC64",x"DCEB",x"C573",x"B5D7",x"BDF7",
									 x"CE79",x"DEFB",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FED7",x"F447",
									 x"EBE2",x"F3E2",x"F442",x"F483",x"F4C3",x"F4E4",x"FD04",x"FD24",x"FD44",x"FD64",
									 x"FD64",x"FD86",x"FE2C",x"FED3",x"FF58",x"FF9A",x"FF9A",x"FF9A",x"FF99",x"FF99",
									 x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAB",x"FE8A",x"FE89",
									 x"FE68",x"FE47",x"FE47",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEA5",x"FEC5",x"FEE5",x"FF05",
									 x"E5C4",x"9321",x"69A1",x"50E0",x"5940",x"61A0",x"6180",x"5920",x"7A86",x"BD32",
									 x"D699",x"F79D",x"F7DE",x"F7DE",x"F7DF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"CE17",x"6AE9",x"4182",
									 x"4160",x"59C0",x"6A41",x"7A81",x"82A1",x"9301",x"9B41",x"A362",x"B382",x"BBA2",
									 x"C3C3",x"C3E3",x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC23",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C423",x"BC23",
									 x"BC02",x"B3E3",x"ABA3",x"9B61",x"B483",x"CDA4",x"EF26",x"FFC7",x"FF86",x"FF46",
									 x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FE85",
									 x"FE65",x"FE45",x"FE04",x"FE05",x"FDE4",x"FDA4",x"FD63",x"FD44",x"F4E3",x"F4A3",
									 x"F462",x"EC64",x"DCEC",x"C593",x"B5D7",x"BDF7",x"CE79",x"DEFB",x"F79E",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FEF7",x"F447",x"EBE2",x"F3E2",x"F442",x"F483",
									 x"F4C3",x"F4E4",x"FD04",x"FD24",x"FD44",x"FD64",x"FD64",x"FDA6",x"FE2C",x"FED3",
									 x"FF58",x"FF9A",x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",
									 x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAB",x"FE8A",x"FE89",x"FE68",x"FE47",x"FE47",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FEA5",x"FEA5",x"FEA5",x"FEC5",x"FEE5",x"FF05",x"E5C4",x"9321",x"69A1",x"50E0",
									 x"5920",x"6180",x"6180",x"5940",x"7A86",x"BD32",x"D699",x"F79D",x"F7DE",x"F7DE",
									 x"F7DF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFDE",x"CE17",x"6AE9",x"41A2",x"4160",x"59E0",x"6A41",x"7A81",
									 x"82A1",x"9301",x"9B41",x"AB62",x"B382",x"BBA2",x"C3C3",x"C3E3",x"C403",x"C403",
									 x"CC23",x"CC23",x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"C443",x"C443",x"C443",x"BC23",x"BC02",x"B3E3",x"ABA3",x"9B62",
									 x"B483",x"CDA4",x"EF26",x"FFC7",x"FF86",x"FF46",x"FF05",x"FEE5",x"FEE5",x"FEE5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE25",x"FE24",x"FE05",
									 x"FDE4",x"FDA4",x"FD84",x"FD44",x"F4E3",x"F4A3",x"F482",x"EC64",x"DCEC",x"C593",
									 x"B5D7",x"BDF7",x"CE59",x"DEFB",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FEF7",x"F447",x"EBE2",x"F3E2",x"F442",x"F483",x"F4C3",x"F4E4",x"FD04",x"FD24",
									 x"FD44",x"FD64",x"FD84",x"FDA6",x"FE2C",x"FED3",x"FF58",x"FF9A",x"FF9A",x"FF9A",
									 x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAB",
									 x"FE8A",x"FE89",x"FE68",x"FE47",x"FE47",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEA5",x"FEC5",
									 x"FEE5",x"FF05",x"E5C4",x"9321",x"69A1",x"50E0",x"5940",x"6180",x"6180",x"6140",
									 x"7A86",x"BD32",x"D699",x"F79D",x"F7DE",x"F7DE",x"F7DF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"CE17",
									 x"6AE9",x"41A2",x"4160",x"59E0",x"6A41",x"7A81",x"82A1",x"9301",x"9B41",x"AB62",
									 x"B382",x"BBA2",x"C3C3",x"C3E3",x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC23",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",
									 x"C443",x"BC23",x"BC02",x"B3E3",x"ABA3",x"9B61",x"B483",x"CDC4",x"EF26",x"FFC7",
									 x"FF86",x"FF46",x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FE85",x"FE85",x"FE65",x"FE25",x"FE24",x"FE05",x"FDE4",x"FDA4",x"FD84",x"FD44",
									 x"F4E3",x"F4A3",x"F482",x"EC84",x"DCEC",x"C593",x"B5D7",x"BDF7",x"CE59",x"DEFB",
									 x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FEF7",x"F447",x"EBE2",x"F3E2",
									 x"F442",x"F483",x"F4C3",x"F4E4",x"FD04",x"FD24",x"FD44",x"FD64",x"FD84",x"FDA6",
									 x"FE2C",x"FED3",x"FF58",x"FF9A",x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",
									 x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAB",x"FE8B",x"FE89",x"FE68",x"FE47",
									 x"FE47",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEA5",x"FEC5",x"FEE5",x"FF05",x"DDC4",x"9321",
									 x"69A1",x"50E0",x"5940",x"6180",x"6180",x"6160",x"7AA7",x"BD52",x"D699",x"F79D",
									 x"F7DE",x"F7DE",x"F7DF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"CE17",x"6AE9",x"4182",x"4160",x"59C0",
									 x"6A41",x"7A81",x"82A1",x"9301",x"9B41",x"AB62",x"B382",x"BBA2",x"C3C2",x"C3E3",
									 x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C443",x"BC23",x"BC02",x"B3E3",
									 x"AB83",x"9B61",x"B483",x"CDC4",x"EF26",x"FFC7",x"FF86",x"FF46",x"FF05",x"FEE5",
									 x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE25",
									 x"FE24",x"FE05",x"FDE4",x"FDA4",x"FD84",x"FD44",x"F4E3",x"F4A3",x"F482",x"EC64",
									 x"DCEC",x"C593",x"B5D7",x"BDF7",x"CE79",x"E71C",x"F79E",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FED7",x"EC67",x"F3E2",x"EC03",x"F442",x"F483",x"F4C3",x"FCE4",
									 x"FD04",x"FD24",x"FD64",x"FD64",x"FD84",x"F5A6",x"FE2B",x"FED2",x"FF58",x"FF9A",
									 x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",
									 x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",
									 x"FEAC",x"FEAC",x"FE8B",x"FE89",x"FE68",x"FE47",x"FE47",x"FE47",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FEA5",x"FEC5",x"FEE5",x"FEE5",x"DDA5",x"9321",x"69A1",x"50E0",x"5940",x"6180",
									 x"6160",x"6160",x"82C6",x"BD72",x"D699",x"F79D",x"F7BE",x"F7DE",x"F7DF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDE",x"C617",x"6AE9",x"4182",x"4160",x"59E0",x"6A41",x"7281",x"82A1",x"9302",
									 x"9B41",x"A362",x"B382",x"BBA2",x"C3C2",x"C3E2",x"C403",x"C403",x"CC23",x"CC23",
									 x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"C443",x"C443",x"C443",x"BC23",x"B402",x"B3C3",x"AB83",x"9B61",x"B483",x"CDC5",
									 x"F746",x"FFC6",x"FF86",x"FF46",x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE24",x"FE24",x"FDE5",x"FDC4",x"FDA4",
									 x"FD63",x"FD23",x"F4E3",x"F4A3",x"F462",x"EC64",x"DCCB",x"C593",x"BDD7",x"BDF8",
									 x"CE79",x"DEFB",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FED7",x"EC68",
									 x"F3E3",x"EC03",x"F442",x"F483",x"F4C3",x"FCE4",x"FD04",x"FD24",x"FD64",x"FD64",
									 x"FD64",x"F5A6",x"FE2B",x"FED2",x"FF58",x"FF9A",x"FF9A",x"FF9A",x"FF99",x"FF99",
									 x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",
									 x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FEAC",x"FE8B",x"FE89",
									 x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEC5",x"FEC4",x"FEC5",
									 x"DDA5",x"9321",x"69A1",x"50E0",x"6140",x"6181",x"6160",x"6180",x"82E7",x"BD73",
									 x"D699",x"F77D",x"F7BE",x"F7DE",x"F7DF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"C5F7",x"62C8",x"4182",
									 x"4180",x"59E0",x"6A62",x"7A81",x"82A1",x"9302",x"9B41",x"A362",x"B382",x"BBA2",
									 x"C3C2",x"C3E2",x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC23",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C423",x"BC23",
									 x"B402",x"B3C3",x"AB82",x"9B60",x"B4A3",x"CDE5",x"F746",x"FFC6",x"FF86",x"FF46",
									 x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FE85",
									 x"FE45",x"FE24",x"FE04",x"FDE5",x"FDC4",x"FDA4",x"FD63",x"FD23",x"F4E3",x"F4A3",
									 x"F462",x"EC65",x"DCCB",x"C573",x"BDD7",x"BDF8",x"CE79",x"DEFB",x"F79E",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FED8",x"EC88",x"F3E3",x"EC03",x"F442",x"F483",
									 x"F4C3",x"FCE4",x"FD04",x"FD24",x"FD44",x"FD64",x"F564",x"F5A6",x"FE2B",x"FED2",
									 x"FF38",x"FF9A",x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",
									 x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FE8C",x"FEAC",x"FEAC",x"FE8B",x"FE89",x"FE68",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FEA5",x"FEC5",x"FEC5",x"FEE6",x"DDA5",x"9301",x"69A1",x"50E0",
									 x"5940",x"6181",x"6160",x"6180",x"8307",x"C573",x"DE99",x"F79D",x"F7BE",x"F7DE",
									 x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFDE",x"C5D6",x"6288",x"4181",x"4180",x"59E0",x"6A62",x"7A81",
									 x"82C2",x"9322",x"9B41",x"A362",x"B382",x"BBA2",x"C3C2",x"C3E2",x"C403",x"C403",
									 x"CC23",x"CC23",x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"CC43",x"C443",x"C443",x"C443",x"C423",x"BC23",x"B402",x"B3C3",x"AB62",x"9B40",
									 x"B4C3",x"D605",x"F746",x"FFC6",x"FF86",x"FF26",x"FF05",x"FEE5",x"FEE5",x"FEE5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE45",x"FE24",x"FE04",x"FDE5",
									 x"FDC4",x"FD84",x"FD63",x"F503",x"F4E3",x"F4A3",x"F463",x"EC65",x"D4CC",x"C573",
									 x"BDD7",x"C618",x"CE79",x"DEFB",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FED8",x"ECA9",x"F404",x"EC03",x"F442",x"F483",x"F4C3",x"FCE3",x"FD04",x"FD24",
									 x"FD44",x"FD64",x"FD64",x"FD86",x"FE2A",x"FEB1",x"FF37",x"FF9A",x"FF9A",x"FF9A",
									 x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF55",x"FF35",x"FF54",
									 x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FEAC",
									 x"FE8B",x"FE89",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEC5",
									 x"FEC5",x"FEC6",x"DDA5",x"8AE1",x"69A1",x"50E0",x"5940",x"6160",x"6160",x"6180",
									 x"8B28",x"C593",x"DEBA",x"F79D",x"F7BE",x"F7DE",x"F7BE",x"FFDF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFBE",x"BDB6",
									 x"5A67",x"4181",x"4180",x"59E0",x"6A61",x"7A81",x"82C1",x"9302",x"9B41",x"A362",
									 x"B382",x"BBA2",x"C3C2",x"C3E2",x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC23",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",
									 x"C423",x"BC23",x"B402",x"B3C3",x"A362",x"9B60",x"BCC3",x"D625",x"F766",x"FFC6",
									 x"FF86",x"FF26",x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FE85",x"FE85",x"FE45",x"FE24",x"FE04",x"FDE5",x"FDC4",x"FDA4",x"FD63",x"FD23",
									 x"F4E3",x"F4A3",x"F483",x"EC86",x"D4EC",x"C574",x"BDD7",x"BE18",x"CE79",x"E71C",
									 x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FEF9",x"F4AA",x"F404",x"EC04",
									 x"F422",x"FC83",x"F4C3",x"F4E3",x"FD04",x"FD24",x"FD44",x"FD64",x"FD64",x"FD85",
									 x"FE2A",x"FEB1",x"FF37",x"FF9A",x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",
									 x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF55",x"FF55",x"FF55",x"FF35",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FEAC",x"FE8B",x"FE89",x"FE68",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEC5",x"FEC5",x"FEC6",x"D584",x"8AC0",
									 x"6181",x"50E0",x"6140",x"6160",x"6160",x"61A0",x"8B48",x"C5B3",x"DEBA",x"F79D",
									 x"F7BE",x"F7BE",x"F7BE",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",
									 x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFBE",x"BD95",x"5A46",x"4181",x"4980",x"5A00",
									 x"6A61",x"7AA1",x"82C1",x"9302",x"9B41",x"A362",x"B382",x"BBA2",x"C3C2",x"C3E2",
									 x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C423",x"BC23",x"B402",x"B3C3",
									 x"A362",x"9B60",x"BD04",x"DE65",x"F786",x"FFC6",x"FF86",x"FF26",x"FF05",x"FEE5",
									 x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE45",x"FE24",
									 x"FE04",x"FDE5",x"FDC4",x"FDA4",x"FD63",x"FD23",x"F4E3",x"F4A3",x"F483",x"EC86",
									 x"D4ED",x"C574",x"BDD7",x"C618",x"D69A",x"E71C",x"F79E",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FF19",x"F4CA",x"F424",x"EC04",x"F422",x"FC83",x"F4A3",x"F4C3",
									 x"F504",x"FD24",x"FD44",x"FD64",x"FD65",x"FD85",x"FE09",x"FEB0",x"FF37",x"FF9A",
									 x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF55",
									 x"FF35",x"FF54",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",
									 x"FEAC",x"FEAC",x"FE8B",x"FE89",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FEA5",x"FEC5",x"FEC5",x"FEA5",x"D544",x"82C0",x"6181",x"50E0",x"6140",x"6160",
									 x"6160",x"61A0",x"8B48",x"C5B3",x"DEBA",x"F79D",x"F7BE",x"F7BE",x"F7BE",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDE",x"FFDF",x"FFFF",x"FFFF",
									 x"FFBE",x"B575",x"5226",x"4161",x"49A0",x"5A00",x"6A61",x"7AA1",x"82C1",x"9302",
									 x"9B41",x"AB62",x"B382",x"BBC2",x"C3E2",x"C3E2",x"C403",x"C403",x"CC23",x"CC23",
									 x"CC23",x"CC23",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"C443",x"C443",x"C422",x"BC02",x"B402",x"B3C3",x"A342",x"9B40",x"C524",x"E6A6",
									 x"FFA7",x"FFA6",x"FF66",x"FF26",x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE45",x"FE24",x"FE04",x"FDE5",x"FDC4",x"FDA4",
									 x"FD63",x"FD23",x"F4E3",x"F4A3",x"F483",x"E487",x"D4ED",x"C594",x"BDD8",x"C618",
									 x"D69A",x"E71C",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF19",x"F4EB",
									 x"F425",x"EC04",x"F422",x"F463",x"F4A3",x"F4E3",x"FD04",x"FD24",x"FD44",x"FD64",
									 x"FD64",x"FD85",x"FDE9",x"FE8F",x"FF37",x"FF7A",x"FF9A",x"FF9A",x"FF99",x"FF99",
									 x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FE8C",x"FE8B",x"FE89",
									 x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FE85",x"FEA5",x"FEC5",x"FEC5",x"FE85",
									 x"D524",x"8281",x"6161",x"50E0",x"6140",x"6160",x"6140",x"61A0",x"8B68",x"C5B3",
									 x"DEBA",x"F77D",x"F79E",x"F7BE",x"F7BF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDE",x"FFDE",x"FFFF",x"FFFF",x"FFDE",x"B574",x"49E5",x"4160",
									 x"49A0",x"5A00",x"6A61",x"7AA1",x"82C1",x"9322",x"A341",x"AB62",x"B382",x"BBC2",
									 x"BBC2",x"C3E2",x"C3E2",x"C403",x"CC23",x"CC23",x"CC23",x"C423",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C443",x"C443",x"C422",x"BC03",
									 x"B3E3",x"B3C2",x"A322",x"9B41",x"C564",x"E706",x"FFA7",x"FFA7",x"FF46",x"FF26",
									 x"FF05",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",
									 x"FE45",x"FE25",x"FE04",x"FDE5",x"FDC4",x"FDA4",x"FD63",x"FD23",x"F4C3",x"F4A3",
									 x"EC64",x"E488",x"CCEE",x"BD94",x"BDD7",x"C618",x"D69A",x"E73C",x"F79E",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF1A",x"F52C",x"F467",x"EC04",x"F422",x"F463",
									 x"F4A3",x"F4E3",x"FD04",x"F504",x"FD44",x"FD65",x"FD84",x"FD85",x"FDE8",x"FE6F",
									 x"FF36",x"FF7A",x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",
									 x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",
									 x"FEAC",x"FE8C",x"FEAC",x"FE8C",x"FE8B",x"FE69",x"FE68",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FEA5",x"FE85",x"FEA5",x"FEC5",x"FEC5",x"FE85",x"D524",x"8281",x"6161",x"5100",
									 x"6140",x"6961",x"6140",x"61C0",x"8B68",x"C5B3",x"DEBA",x"F77D",x"F79E",x"F79E",
									 x"F7BF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDE",x"FFDF",
									 x"FFFF",x"FFFF",x"FFBE",x"B574",x"49C4",x"3960",x"49A0",x"5A00",x"6A61",x"7AA1",
									 x"82C1",x"9302",x"A341",x"AB62",x"B382",x"BBC2",x"BBC2",x"C3E2",x"C3E2",x"C403",
									 x"CC23",x"CC23",x"C423",x"C423",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",
									 x"C443",x"C443",x"C443",x"C442",x"BC22",x"BC03",x"B3E3",x"ABC2",x"A342",x"9B41",
									 x"CD84",x"EF46",x"FFC7",x"FFA7",x"FF46",x"FF26",x"FEE5",x"FEE5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE45",x"FE25",x"FE05",x"FDE5",
									 x"FDC4",x"F583",x"FD64",x"FD03",x"F4C3",x"F4A3",x"EC84",x"E489",x"CD0E",x"BD93",
									 x"BDD7",x"C638",x"D6BA",x"E73C",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FF1A",x"F54D",x"F488",x"EC25",x"F422",x"F463",x"F4A3",x"F4E3",x"FD04",x"F504",
									 x"FD44",x"FD64",x"FD85",x"FD85",x"FDC7",x"FE6E",x"FF36",x"FF7A",x"FF9A",x"FF9A",
									 x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FE8C",
									 x"FE8B",x"FE69",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FE85",x"FEA5",x"FEC5",
									 x"FEC5",x"FE85",x"D524",x"8261",x"6161",x"5100",x"6140",x"6961",x"6140",x"61C0",
									 x"8368",x"C593",x"DEBA",x"EF7D",x"F79E",x"F79E",x"F7BE",x"F7DF",x"FFDF",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDE",x"FFDF",x"FFFF",x"FFFF",x"FFBE",x"B553",
									 x"41C4",x"4160",x"49C0",x"5A00",x"6A61",x"7AA1",x"82C1",x"9322",x"A341",x"AB62",
									 x"B382",x"BBC2",x"BBC2",x"C3E2",x"C3E2",x"C403",x"CC23",x"CC23",x"C423",x"C423",
									 x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C443",x"C443",x"C442",
									 x"BC22",x"BC03",x"ABE3",x"ABC2",x"9B42",x"9B61",x"CDC5",x"EF46",x"FFC7",x"FFA6",
									 x"FF26",x"FF06",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",
									 x"FE85",x"FE65",x"FE45",x"FE25",x"FE04",x"FDC4",x"FDA4",x"F583",x"F563",x"FD04",
									 x"F4C3",x"ECA3",x"EC85",x"E4A9",x"CD0F",x"BD94",x"BDF7",x"C659",x"D6BA",x"EF5D",
									 x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF5B",x"F58F",x"F4A9",x"EC26",
									 x"F423",x"F463",x"F4A3",x"F4E3",x"FD04",x"F504",x"FD44",x"FD64",x"FD65",x"FD84",
									 x"FDA6",x"FE4C",x"FF15",x"FF7A",x"FF9A",x"FF9A",x"FF99",x"FF99",x"FF99",x"FF99",
									 x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FEAD",x"FEAD",x"FEAD",
									 x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FE8C",x"FE8B",x"FE69",x"FE68",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FEA5",x"FEA5",x"FE85",x"FEA5",x"FEC5",x"FEC5",x"F685",x"CD03",x"8261",
									 x"6161",x"5100",x"6140",x"6961",x"6140",x"61C0",x"8B68",x"C593",x"D6BA",x"EF7D",
									 x"F79D",x"F79E",x"F7BE",x"F7BF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"F7DE",
									 x"FFDE",x"FFDF",x"FFFF",x"FFFF",x"F7BD",x"AD33",x"41A4",x"4160",x"49C0",x"5A00",
									 x"6A61",x"7AA1",x"82C2",x"9322",x"A341",x"AB62",x"B382",x"BBC2",x"BBC2",x"C3E2",
									 x"C3E3",x"C403",x"CC23",x"CC23",x"CC23",x"C423",x"CC43",x"CC43",x"CC43",x"CC43",
									 x"CC43",x"C443",x"C443",x"C443",x"C422",x"C422",x"C422",x"B3E3",x"ABC3",x"ABA2",
									 x"9B41",x"A3C1",x"D605",x"F787",x"FFC7",x"FF86",x"FF26",x"FF06",x"FEE5",x"FEE5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE05",
									 x"FE04",x"FDC4",x"FDA4",x"FD83",x"FD44",x"F504",x"F4A3",x"F4A4",x"EC86",x"E4CA",
									 x"CD2F",x"BD94",x"BDF8",x"CE59",x"DEDB",x"EF5D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"F77C",x"F5B0",x"F4CA",x"EC47",x"F423",x"F443",x"F4A3",x"F4C3",
									 x"FD04",x"F504",x"FD44",x"FD64",x"FD65",x"FD64",x"FD85",x"FE2B",x"FF14",x"FF7A",
									 x"FF9A",x"FF9A",x"FF99",x"FF79",x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",
									 x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FEF0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FE8C",
									 x"FEAC",x"FE8C",x"FE8B",x"FE69",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FE85",
									 x"FEA5",x"FEC5",x"FEC5",x"F664",x"CCE3",x"8260",x"6161",x"5100",x"6140",x"6961",
									 x"6140",x"61C0",x"8B88",x"C5B3",x"D6BA",x"EF7D",x"EF7D",x"F79E",x"F7BE",x"F7BF",
									 x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"FFDE",x"FFDF",x"FFFF",
									 x"F79D",x"AD13",x"3983",x"4160",x"49C0",x"5A20",x"7282",x"7AA1",x"82C2",x"9322",
									 x"A341",x"AB62",x"B382",x"BBA2",x"BBC2",x"C3E2",x"C3E3",x"C403",x"CC23",x"CC23",
									 x"CC23",x"C423",x"CC43",x"CC43",x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C443",
									 x"C443",x"BC22",x"BC22",x"B3E3",x"ABC3",x"A381",x"9B62",x"A402",x"D645",x"F7A7",
									 x"FFC6",x"FF86",x"FF26",x"FF06",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE05",x"FDE4",x"FDC4",x"FDA4",x"FD84",
									 x"FD44",x"FCE4",x"F4A4",x"F4A4",x"EC86",x"DCCB",x"CD30",x"BD94",x"BDF8",x"CE79",
									 x"DEDB",x"EF5D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F77C",x"FDD1",
									 x"F4EB",x"EC47",x"F403",x"F443",x"F4A3",x"F4C3",x"FD04",x"F504",x"FD44",x"FD64",
									 x"FD65",x"FD64",x"FD64",x"F60A",x"FEF3",x"FF79",x"FF9A",x"FF9A",x"FF99",x"FF79",
									 x"FF99",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FEF0",x"FECF",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FEAD",
									 x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAC",x"FE8C",x"FE8B",x"FE69",
									 x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FE85",x"FEA5",x"FEC5",x"FEC5",x"F664",
									 x"CCE3",x"8240",x"6161",x"5100",x"6140",x"6960",x"6140",x"61C0",x"8B88",x"C5B3",
									 x"DEBA",x"EF5D",x"EF7D",x"F79E",x"F79E",x"F7BF",x"F7BE",x"F7BE",x"F7BE",x"F7BE",
									 x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"FFDF",x"FFFF",x"F79D",x"A4F2",x"3943",x"4160",
									 x"51E0",x"6220",x"7282",x"7AA1",x"82C2",x"9322",x"A341",x"AB62",x"B382",x"BBA2",
									 x"BBC2",x"C3E2",x"C3E3",x"C403",x"CC23",x"CC23",x"CC23",x"C423",x"CC43",x"CC43",
									 x"CC43",x"CC43",x"CC43",x"C443",x"C443",x"C443",x"C422",x"BC22",x"BC22",x"B3E2",
									 x"ABA3",x"A381",x"A382",x"AC63",x"DE85",x"FFA7",x"FFA6",x"FF65",x"FF26",x"FF06",
									 x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",
									 x"FE45",x"FE05",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD44",x"FCE4",x"F4A4",x"F4A4",
									 x"ECA7",x"DCEC",x"CD51",x"BD95",x"BE18",x"CE9A",x"DEFB",x"EF7D",x"FFDF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF7B",x"F613",x"F50D",x"EC67",x"F423",x"F462",
									 x"F482",x"FCC3",x"FCE4",x"FD04",x"FD24",x"FD44",x"FD85",x"FD64",x"FD85",x"FE09",
									 x"FED1",x"FF58",x"FF9A",x"FF9A",x"FF79",x"FF79",x"FF99",x"FF99",x"FF99",x"FF99",
									 x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF35",x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FEAD",x"FEAD",x"FEAD",x"FE8C",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAB",x"FE8B",x"FE6A",x"FE68",x"FE67",x"FE46",x"FE46",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FEA5",x"FEA5",x"FEA4",x"FEE5",x"FEC5",x"F664",x"C4C3",x"7A60",x"6161",x"5920",
									 x"6140",x"6141",x"6140",x"61C1",x"8B89",x"C5D3",x"DEBA",x"EF7D",x"EF7D",x"EF7D",
									 x"F79E",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",
									 x"F7DF",x"FFDF",x"F77D",x"A4D2",x"3122",x"3961",x"51E0",x"6220",x"7281",x"7AA1",
									 x"8AC2",x"9B22",x"A341",x"AB62",x"B382",x"BBC2",x"BBE2",x"C3E3",x"C403",x"C403",
									 x"CC23",x"CC23",x"CC23",x"CC23",x"CC23",x"CC43",x"CC42",x"CC42",x"CC42",x"C443",
									 x"C443",x"C443",x"C423",x"BC23",x"BC02",x"B402",x"ABA2",x"A362",x"A3A2",x"BCE3",
									 x"E6C6",x"FFA7",x"FFA7",x"FF45",x"FF05",x"FF06",x"FEE5",x"FEE5",x"FEC5",x"FEC5",
									 x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE65",x"FE45",x"FE25",x"FDE5",x"FDC4",
									 x"FDA4",x"FD64",x"FD24",x"F4E4",x"F4A4",x"F484",x"E4A8",x"DD0D",x"CD51",x"BD95",
									 x"BE19",x"D69A",x"E71C",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FF9C",x"F675",x"F54F",x"F488",x"EC24",x"F462",x"F462",x"F4A3",x"FCC3",x"FD04",
									 x"FD24",x"FD44",x"FD65",x"FD85",x"FD85",x"FDE8",x"FEAF",x"FF37",x"FF9A",x"FF9A",
									 x"FF79",x"FF79",x"FF79",x"FF99",x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",
									 x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FE8A",x"FE69",x"FE67",x"FE66",x"FE66",x"FE47",x"FE67",x"FE67",x"FE67",
									 x"FE67",x"FE67",x"FE67",x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",
									 x"FE67",x"FE66",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEA4",x"FEE5",
									 x"F6C5",x"EE64",x"BC83",x"7A40",x"6140",x"5920",x"6160",x"6141",x"6140",x"69C1",
									 x"93CA",x"C5D4",x"DEDB",x"EF7D",x"EF7D",x"F79E",x"F79E",x"F7BE",x"F7BE",x"F7BE",
									 x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"FFBE",x"F7BE",x"FFFF",x"F7DE",x"E71B",x"9C70",
									 x"3102",x"3960",x"51E0",x"6220",x"7A81",x"7AC1",x"8AE2",x"9B22",x"A341",x"AB62",
									 x"B382",x"BBC2",x"C3E2",x"C3E3",x"C403",x"C403",x"C403",x"CC23",x"CC23",x"CC23",
									 x"CC22",x"CC22",x"C442",x"C442",x"C442",x"C443",x"C443",x"C443",x"C443",x"BC23",
									 x"BC03",x"B3E2",x"AB82",x"9B22",x"A3C2",x"CD84",x"EF06",x"FFA7",x"FFA7",x"FF45",
									 x"FF05",x"FF05",x"FEE6",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",
									 x"FE65",x"FE45",x"FE45",x"FE05",x"FDE4",x"FDA4",x"FD84",x"FD64",x"FD24",x"F4E4",
									 x"F4A4",x"F484",x"E4C9",x"D52E",x"CD72",x"BDB5",x"C639",x"D6BB",x"E71C",x"F79E",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"FEB7",x"F590",x"F4A9",
									 x"EC24",x"F442",x"F442",x"F4A3",x"FCC4",x"FD04",x"FD24",x"FD44",x"FD64",x"FD85",
									 x"FD85",x"FDE8",x"FE8E",x"FF16",x"FF99",x"FF9A",x"FF79",x"FF79",x"FF79",x"FF99",
									 x"FF99",x"FF99",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FECD",x"FECB",x"FEAA",x"FEA8",
									 x"FEC8",x"FEC8",x"FEC8",x"FEC8",x"FEC8",x"FEA8",x"FEA8",x"FE87",x"FE67",x"FE67",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE66",x"FE67",x"FE47",
									 x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEA4",x"FEE5",x"FEC5",x"E644",x"B462",x"7200",
									 x"5920",x"5920",x"6160",x"6140",x"6140",x"69E2",x"9BEB",x"CDF5",x"DEDB",x"EF5D",
									 x"EF7D",x"F79E",x"F79E",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",
									 x"F7BE",x"F7BE",x"F7DF",x"F7BE",x"DEB9",x"942F",x"3102",x"4160",x"51E0",x"6220",
									 x"7A81",x"82C1",x"8AE1",x"9B22",x"A361",x"AB62",x"B382",x"BBC2",x"C3E2",x"C3E3",
									 x"C403",x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC22",x"CC22",x"C442",x"C442",
									 x"C442",x"C443",x"C443",x"C443",x"C423",x"BC02",x"B402",x"B3E2",x"A382",x"9301",
									 x"A3C2",x"D605",x"F746",x"FFC7",x"FF86",x"FF46",x"FF05",x"FF06",x"FEE6",x"FEC5",
									 x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE45",x"FE25",x"FE05",
									 x"FDE4",x"FDA4",x"FD84",x"FD44",x"FD23",x"F4C3",x"F4A4",x"F485",x"DCCA",x"D550",
									 x"CD93",x"BDB6",x"C659",x"DEDB",x"E73C",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFBD",x"F6F9",x"F5D2",x"F4CB",x"EC25",x"F442",x"F462",x"FCA3",
									 x"FCC4",x"FD04",x"FD24",x"FD44",x"FD64",x"FD84",x"FD85",x"FDE7",x"FE8D",x"FF15",
									 x"FF99",x"FF9A",x"FF79",x"FF79",x"FF79",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF55",
									 x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECE",x"FEAE",x"FECD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FECC",x"FECC",x"FECC",x"FECB",x"FEA9",x"FEA9",x"FEA8",x"F6C8",x"F6C8",x"FEC8",
									 x"FEC8",x"FEC8",x"FEC8",x"FEA7",x"FE87",x"FEA8",x"FE88",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE67",x"FE67",x"FE66",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",
									 x"FEA4",x"FEE5",x"FEC5",x"E624",x"B423",x"69E1",x"5900",x"5900",x"6160",x"6141",
									 x"6120",x"69E3",x"9C2C",x"CE16",x"DEDB",x"EF5D",x"EF7D",x"EF7D",x"F79E",x"F79E",
									 x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7DF",x"EF9D",
									 x"D678",x"8C0E",x"3102",x"4181",x"59E0",x"6220",x"7A81",x"82C1",x"8AE2",x"9B22",
									 x"AB61",x"B362",x"BB82",x"BBC2",x"C3E2",x"C3E3",x"C403",x"C403",x"C403",x"CC23",
									 x"CC23",x"CC23",x"CC22",x"CC22",x"C442",x"C442",x"C442",x"C443",x"C443",x"C443",
									 x"C423",x"BC02",x"B3E3",x"B3E3",x"A362",x"9300",x"A3E2",x"DE66",x"F786",x"FFC7",
									 x"FF86",x"FF26",x"FF05",x"FEE6",x"FEE6",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",
									 x"FEA5",x"FE85",x"FE65",x"FE45",x"FE25",x"FE05",x"FDE4",x"FDA4",x"FD84",x"FD44",
									 x"FD24",x"F4C3",x"F484",x"EC86",x"DCCB",x"CD71",x"C5B4",x"BDD6",x"CE59",x"DEFB",
									 x"EF5D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",x"FF3A",
									 x"F634",x"F50C",x"EC25",x"F422",x"F442",x"FC83",x"FCC4",x"FD04",x"FD24",x"FD44",
									 x"FD64",x"FD64",x"FD84",x"FDE7",x"FE6C",x"FEF4",x"FF99",x"FF9A",x"FF79",x"FF79",
									 x"FF79",x"FF99",x"FF99",x"FF99",x"FF99",x"FF99",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",
									 x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FEAE",x"FEAD",x"FEAD",
									 x"FECD",x"FEAC",x"FECC",x"FECC",x"FEEC",x"FEED",x"FECD",x"F68C",x"EE4B",x"E5EA",
									 x"DDA8",x"D587",x"D587",x"D587",x"D587",x"DDA7",x"E5E7",x"EE28",x"F668",x"FEC9",
									 x"FF0A",x"FF0A",x"FEE9",x"FEA8",x"FE88",x"FE87",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE66",
									 x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA4",x"FEE5",x"F6C5",x"E604",
									 x"ABE3",x"69A1",x"5900",x"5920",x"6160",x"6141",x"5920",x"7224",x"A46E",x"CE37",
									 x"DEFB",x"EF5D",x"EF7D",x"EF7D",x"EF7D",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",
									 x"F79E",x"F79E",x"F79E",x"F7BE",x"F7DF",x"EF5C",x"C616",x"83CD",x"3122",x"4181",
									 x"59E0",x"6A20",x"7A81",x"82C1",x"8AE2",x"9B22",x"AB61",x"B382",x"BB82",x"BBC2",
									 x"C3E2",x"C3E3",x"C403",x"C403",x"C403",x"CC23",x"CC23",x"CC23",x"CC22",x"CC22",
									 x"C442",x"C442",x"C442",x"C442",x"C443",x"C443",x"BC23",x"BC02",x"BC03",x"B3C3",
									 x"A362",x"9300",x"AC42",x"EEE7",x"F7A6",x"FFC6",x"FF86",x"FF26",x"FEE6",x"FEE6",
									 x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE45",
									 x"FE25",x"FE05",x"FDC4",x"FDA4",x"FD84",x"FD43",x"FD04",x"FCC3",x"FC84",x"EC86",
									 x"D4EC",x"CD93",x"C5D6",x"C5F7",x"CE79",x"DEFB",x"EF5D",x"FFDF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF9C",x"FE76",x"F54E",x"EC46",x"F402",
									 x"F442",x"F483",x"FCC3",x"FCE4",x"FD24",x"FD44",x"FD64",x"FD64",x"FD84",x"FDC6",
									 x"F62B",x"FED3",x"FF99",x"FF9A",x"FF79",x"FF79",x"FF79",x"FF99",x"FF99",x"FF99",
									 x"FF99",x"FF99",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FEAE",x"FECE",x"FEAE",x"FEAD",x"FEAD",x"FECD",x"FEED",x"FEED",x"FEED",
									 x"F6AC",x"E62B",x"D589",x"C508",x"B486",x"A405",x"9BA4",x"9363",x"9322",x"9342",
									 x"9342",x"9B82",x"ABE4",x"B465",x"BCE5",x"D5A7",x"DE28",x"E688",x"FF09",x"FF09",
									 x"FEE9",x"FEA8",x"FE87",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE66",x"FE67",x"FE47",x"FE47",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FEA5",x"FEA4",x"FEE5",x"F6C4",x"DDC4",x"A3C3",x"6160",x"58E0",x"5920",
									 x"6180",x"6140",x"5900",x"7224",x"ACAF",x"D678",x"DEFB",x"EF5D",x"EF5D",x"EF7D",
									 x"EF7D",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"F7BE",
									 x"F7DF",x"E71B",x"B574",x"7B6B",x"3121",x"49A1",x"59E0",x"6A20",x"7A81",x"82C1",
									 x"92E2",x"A322",x"AB61",x"B382",x"BB83",x"BBC2",x"C3E2",x"C3E3",x"C403",x"C403",
									 x"C403",x"CC23",x"CC23",x"CC23",x"CC22",x"CC22",x"C442",x"C442",x"C442",x"C422",
									 x"C443",x"C423",x"BC23",x"BC02",x"B3E3",x"ABA2",x"A362",x"9B61",x"B4C4",x"F768",
									 x"F7C6",x"FFC6",x"FF66",x"FF06",x"FEE6",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",
									 x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE45",x"FE25",x"FDE4",x"FDC4",x"FDA4",
									 x"FD63",x"FD43",x"FD03",x"FCA3",x"FC84",x"ECA7",x"D50D",x"C593",x"C5D6",x"C617",
									 x"D699",x"E71C",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FF9D",x"FEB8",x"F5B0",x"EC67",x"F403",x"F422",x"F483",x"FCC3",x"FCE3",
									 x"FD04",x"FD24",x"FD45",x"FD64",x"FD85",x"FDA6",x"F608",x"FEB1",x"FF79",x"FF9B",
									 x"FF7A",x"FF99",x"FF99",x"FF7A",x"FF79",x"FF99",x"FF99",x"FF99",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF54",
									 x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FEAE",x"FECE",
									 x"FECE",x"FEAD",x"FECD",x"FEED",x"FECC",x"F68C",x"DDCA",x"BCC8",x"A3E6",x"9365",
									 x"8303",x"7A82",x"7241",x"61E0",x"61C0",x"69E0",x"69E0",x"7200",x"7A82",x"82E2",
									 x"9363",x"A404",x"B4C5",x"CD66",x"E689",x"F72A",x"FF29",x"FF09",x"FEC7",x"FEA7",
									 x"FE67",x"FE47",x"FE48",x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",
									 x"FE67",x"FE66",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FF06",
									 x"F6C4",x"DDA4",x"A3A3",x"6140",x"58E0",x"6120",x"6961",x"6140",x"5900",x"7245",
									 x"ACD0",x"D698",x"DF1B",x"EF5D",x"EF5D",x"EF7D",x"EF7D",x"EF9E",x"F79E",x"F79E",
									 x"F79E",x"F79E",x"F79E",x"F79E",x"F79D",x"F7BE",x"FFDF",x"DEDA",x"A4F2",x"732A",
									 x"3101",x"49A1",x"5A00",x"6A40",x"7A81",x"82C2",x"9302",x"9B42",x"AB61",x"B382",
									 x"BB83",x"BBC2",x"C3E2",x"C3E3",x"C403",x"C403",x"C403",x"C402",x"CC22",x"CC22",
									 x"CC22",x"CC42",x"C442",x"C442",x"C443",x"C443",x"C422",x"BC22",x"BC22",x"B3E2",
									 x"B3C2",x"AB82",x"A362",x"A3E2",x"C543",x"FF88",x"FFC6",x"FFA6",x"FF45",x"FEE6",
									 x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",
									 x"FE45",x"FE45",x"FE25",x"FDE4",x"FDC4",x"FD84",x"FD64",x"F523",x"FCE3",x"F483",
									 x"F484",x"E4A9",x"D52E",x"BD94",x"BDD7",x"C618",x"D69A",x"E73C",x"EF7D",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FEF9",x"FDF2",
									 x"EC88",x"F403",x"EC22",x"F463",x"FCA3",x"FCE3",x"FD04",x"FD24",x"FD45",x"FD64",
									 x"FD85",x"FDA6",x"F5E7",x"FE8F",x"FF78",x"FF9B",x"FF9B",x"FF9A",x"FF99",x"FF7A",
									 x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF55",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEEE",x"FECD",
									 x"E5EA",x"CD49",x"AC06",x"82E3",x"7241",x"7241",x"6A21",x"6A21",x"6A21",x"6A00",
									 x"6A00",x"7220",x"7220",x"7241",x"7A41",x"7A61",x"7A81",x"7AA1",x"8B03",x"9BA4",
									 x"BCE6",x"DE28",x"F72B",x"FF4B",x"FF2A",x"FEE8",x"FE87",x"FE68",x"FE48",x"FE48",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE66",x"FE67",x"FE47",
									 x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FF06",x"F6C5",x"D5A4",x"9B83",x"5940",
									 x"50E0",x"6141",x"6961",x"6140",x"5100",x"6A46",x"ACF1",x"D699",x"E71C",x"E75C",
									 x"EF5D",x"EF7D",x"EF7D",x"EF9D",x"EF7D",x"EF7D",x"EF7D",x"F79E",x"F79E",x"F79E",
									 x"F79E",x"F7BE",x"FFDF",x"D69A",x"9450",x"6AE8",x"3921",x"49A1",x"5A00",x"6A60",
									 x"7A81",x"82E2",x"9302",x"9B42",x"AB61",x"B382",x"BBA3",x"BBC2",x"C3E2",x"CBE3",
									 x"CC03",x"CC03",x"C402",x"C402",x"CC22",x"CC22",x"CC23",x"C443",x"C443",x"C443",
									 x"C443",x"C443",x"C422",x"BC22",x"BC22",x"B3E2",x"B3E3",x"A342",x"A362",x"B463",
									 x"CDC3",x"FF87",x"FFC7",x"FFA6",x"FF25",x"FEE6",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE44",x"FE25",x"FE05",x"FDE4",
									 x"FDC4",x"FD84",x"FD44",x"F523",x"FCE3",x"F4A3",x"EC85",x"E4CA",x"D54F",x"BD94",
									 x"BDD7",x"C638",x"D6BA",x"E73C",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FF3B",x"FE34",x"ECAA",x"F424",x"F422",x"F463",
									 x"F4A3",x"FCE3",x"FD04",x"FD24",x"FD45",x"FD64",x"FD65",x"FD85",x"F5C6",x"FE4D",
									 x"FF57",x"FF9A",x"FF9A",x"FF9A",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF56",x"FF56",x"FF56",x"FF36",x"FF55",x"FF55",x"FF55",x"FF35",
									 x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FEED",x"FEED",x"F6AD",x"DDCB",x"AC26",x"9345",x"7262",x"59A0",
									 x"5980",x"61A0",x"6A00",x"7240",x"7A81",x"82A2",x"82A2",x"8AC2",x"8AC2",x"8AC1",
									 x"8281",x"8281",x"7A41",x"7221",x"71E1",x"7A21",x"82C2",x"AC65",x"D5C9",x"E68A",
									 x"FF4B",x"FF29",x"FF09",x"FEC8",x"FE88",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",
									 x"FE47",x"FE67",x"FE67",x"FE66",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FEA5",x"FF06",x"F6A4",x"D564",x"9342",x"5900",x"50C0",x"6141",x"6981",x"6140",
									 x"5900",x"7266",x"B512",x"D6B9",x"E73C",x"E73C",x"E75C",x"EF5D",x"EF7D",x"EF7D",
									 x"EF7D",x"EF7D",x"EF7D",x"F79E",x"F79E",x"F79D",x"F79D",x"F79E",x"FFDF",x"D659",
									 x"83ED",x"5A87",x"3941",x"51C1",x"5A00",x"6A60",x"7AA1",x"8AE2",x"9302",x"A342",
									 x"AB81",x"B382",x"BBA3",x"BBC2",x"C3E2",x"CBE3",x"CC03",x"CC03",x"C402",x"C402",
									 x"CC22",x"CC23",x"CC23",x"C423",x"C423",x"C423",x"C423",x"C423",x"BC22",x"BC22",
									 x"B402",x"B3C2",x"ABC3",x"9B00",x"A3A2",x"C525",x"DE65",x"FFA7",x"FFC6",x"FF66",
									 x"FF25",x"FEE6",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",
									 x"FE65",x"FE45",x"FE24",x"FE24",x"FE05",x"FDC4",x"FDA4",x"FD84",x"F544",x"F503",
									 x"FCC3",x"F483",x"ECA6",x"E4EC",x"CD51",x"BDB5",x"BDF7",x"CE58",x"DEDB",x"EF5D",
									 x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",
									 x"FF7C",x"FE75",x"ECEB",x"EC25",x"F423",x"F463",x"F4A3",x"FCC3",x"FD04",x"FD04",
									 x"FD25",x"FD64",x"FD65",x"FD65",x"FDA5",x"FE2C",x"FF15",x"FF79",x"FF7A",x"FF9A",
									 x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF55",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",
									 x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FF12",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FEEF",x"FEEE",x"FECE",x"FECD",x"FEED",x"F68C",
									 x"DDCB",x"AC27",x"7261",x"61C1",x"61A1",x"61C1",x"7201",x"7A41",x"7A61",x"8281",
									 x"82A1",x"82A1",x"8AC1",x"8AC1",x"8AC1",x"92C1",x"92C1",x"92C1",x"8AC1",x"8AA1",
									 x"8AA1",x"8262",x"7A40",x"82C1",x"9BC3",x"BD26",x"EEEA",x"FF6B",x"FF4A",x"FEE9",
									 x"FEA8",x"FE87",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE66",
									 x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA4",x"FF06",x"F6A5",x"CD44",
									 x"8B02",x"50E0",x"50C0",x"6141",x"6981",x"6140",x"5100",x"7287",x"B533",x"D6DA",
									 x"E73C",x"E73C",x"E73C",x"EF5D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",
									 x"EF7D",x"EF7D",x"F79D",x"F79E",x"FFDF",x"CE38",x"7B8C",x"5245",x"4141",x"51C0",
									 x"6220",x"6A40",x"7AA1",x"8AE1",x"9302",x"A342",x"AB81",x"B382",x"BBA3",x"BBC2",
									 x"C3E2",x"CBE3",x"CC03",x"CC03",x"C403",x"C402",x"C423",x"CC23",x"CC23",x"C423",
									 x"C423",x"C423",x"C423",x"C423",x"BC22",x"BC02",x"B403",x"ABC2",x"ABA2",x"92E0",
									 x"A3C2",x"D5C5",x"EEE6",x"FFC7",x"FFA7",x"FF45",x"FF05",x"FEE6",x"FEC6",x"FEC5",
									 x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE44",x"FE24",x"FE24",
									 x"FDE4",x"FDC4",x"FDA4",x"FD64",x"FD43",x"F503",x"FCA2",x"F484",x"ECA7",x"DD0D",
									 x"CD72",x"BDB6",x"BDF8",x"CE59",x"DEFB",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"FED7",x"ED0D",x"EC47",
									 x"F423",x"F443",x"F483",x"F4A3",x"FCE4",x"FD04",x"FD24",x"FD64",x"FD65",x"FD65",
									 x"FD84",x"FE0A",x"FEF3",x"FF78",x"FF7A",x"FF9A",x"FF99",x"FF79",x"FF79",x"FF79",
									 x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",x"FF36",x"FF55",x"FF55",
									 x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FEEF",x"FECE",x"FECE",x"FF0E",x"FECE",x"E5EC",x"BCC9",x"7AC3",x"59A0",x"5980",
									 x"61A0",x"7201",x"7A41",x"8261",x"8281",x"82A1",x"8AC1",x"8AE1",x"92E2",x"92E1",
									 x"92E1",x"92C2",x"92C2",x"92E1",x"92E1",x"92E1",x"92E0",x"8AA0",x"8260",x"8260",
									 x"8AC1",x"9BA3",x"CDE8",x"F74B",x"FF8C",x"FF4A",x"FEC8",x"FEA8",x"FE87",x"FE67",
									 x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE66",x"FE67",x"FE47",x"FE47",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FEA5",x"FEA5",x"FF06",x"EE85",x"C503",x"8AC2",x"50E0",x"50C0",x"6140",
									 x"6980",x"6140",x"5100",x"7287",x"BD54",x"DEDB",x"E73C",x"E73C",x"E73C",x"EF5D",
									 x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"F79E",
									 x"FFDF",x"C617",x"6B0A",x"4A04",x"4160",x"51E0",x"6220",x"6A40",x"82C2",x"8AE1",
									 x"9302",x"A342",x"AB81",x"BBA2",x"BBA2",x"C3C2",x"C3E2",x"CBE3",x"CC03",x"CC03",
									 x"C403",x"C402",x"C423",x"C423",x"CC23",x"C423",x"C443",x"C423",x"C423",x"C423",
									 x"BC23",x"BC03",x"B3E3",x"ABA2",x"A362",x"9320",x"AC42",x"DE46",x"F746",x"FFC7",
									 x"FF86",x"FF25",x"FF06",x"FEE6",x"FEC6",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",
									 x"FE85",x"FE65",x"FE65",x"FE44",x"FE24",x"FE04",x"FDE4",x"FDC4",x"FDA4",x"FD64",
									 x"FD43",x"FCE3",x"F4A3",x"EC84",x"E4C8",x"D52F",x"CD94",x"BDB6",x"BDF8",x"CE59",
									 x"E71C",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFE",x"FF19",x"F56F",x"EC48",x"F403",x"F422",x"F483",x"F4A3",
									 x"FCE4",x"FCE4",x"FD24",x"FD44",x"FD65",x"FD65",x"FDA3",x"FDE9",x"FED2",x"FF77",
									 x"FF9A",x"FF9A",x"FF9A",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",
									 x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",
									 x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FEEF",x"FECE",x"FEEE",x"FEED",
									 x"E64C",x"B488",x"8B25",x"59A0",x"59A0",x"6A01",x"7221",x"7A61",x"8281",x"8AA1",
									 x"8AC1",x"8AC1",x"92E2",x"9302",x"92E2",x"9B02",x"9302",x"9B02",x"9B02",x"9B02",
									 x"9B02",x"9B02",x"9B22",x"9301",x"9301",x"8AA1",x"7A00",x"7A40",x"A404",x"DE6A",
									 x"FF8C",x"FF8B",x"FF09",x"FEC8",x"FE88",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",
									 x"FE67",x"FE66",x"FE67",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FF06",
									 x"EE85",x"C4E3",x"82A1",x"50C0",x"50C0",x"6140",x"6980",x"6140",x"5120",x"7AA8",
									 x"BD75",x"DEDC",x"E73C",x"E73C",x"E73C",x"E75D",x"EF5D",x"EF7D",x"EF5D",x"EF5D",
									 x"EF5D",x"EF7D",x"EF7D",x"EF7D",x"EF7D",x"F79E",x"FFDF",x"BDD6",x"5AA8",x"41A2",
									 x"4160",x"59E0",x"6220",x"7240",x"82C2",x"8AE1",x"9302",x"A342",x"B381",x"BBA2",
									 x"BBA2",x"C3C2",x"C3E2",x"CBE3",x"CC03",x"CC03",x"C403",x"C402",x"C403",x"C423",
									 x"CC23",x"C423",x"C423",x"C423",x"C423",x"C423",x"BC02",x"BC03",x"B3C3",x"A362",
									 x"9B42",x"9B61",x"B4C3",x"E6C6",x"F786",x"FFA6",x"FF66",x"FF06",x"FF06",x"FEE6",
									 x"FEC6",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE44",
									 x"FE24",x"FE04",x"FDE4",x"FDA4",x"FD83",x"FD44",x"F523",x"F4E2",x"F4A2",x"EC85",
									 x"E4E9",x"D550",x"C5B4",x"BDB7",x"C618",x"D699",x"E73C",x"F7BE",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF9C",
									 x"F5F2",x"F469",x"F424",x"F422",x"F462",x"F4A3",x"F4E4",x"F504",x"FD24",x"FD44",
									 x"FD64",x"FD64",x"FD84",x"FDC8",x"FE8F",x"FF76",x"FF7A",x"FF9B",x"FF9A",x"FF79",
									 x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FEEE",x"FECE",x"FEED",x"CD4A",x"7283",x"61C2",x"59A0",
									 x"61E1",x"7221",x"7A41",x"8281",x"8281",x"8AA1",x"92C1",x"92E2",x"92E2",x"9B02",
									 x"9B02",x"9B22",x"9B22",x"A322",x"A322",x"9B22",x"9B22",x"9B02",x"9B02",x"9B22",
									 x"9301",x"92C1",x"8A81",x"7A40",x"82A1",x"BD27",x"DEA9",x"FF8B",x"FF8A",x"FF09",
									 x"FEA8",x"FE67",x"FE47",x"FE67",x"FE47",x"FE67",x"FE67",x"FE66",x"FE67",x"FE47",
									 x"FE47",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",
									 x"FE85",x"FE65",x"FE85",x"FE85",x"FEA5",x"FEE6",x"EE44",x"BCA3",x"8261",x"50C0",
									 x"50C0",x"6160",x"69A0",x"6140",x"5920",x"7AC8",x"BD95",x"DEDB",x"E73C",x"E73C",
									 x"E73C",x"E75D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",
									 x"EF7D",x"F79E",x"FFDF",x"BD95",x"49E5",x"3941",x"4980",x"5A00",x"6240",x"7261",
									 x"82C2",x"9301",x"9B21",x"A342",x"B382",x"BBA2",x"BBA3",x"C3C2",x"C3E2",x"CBE2",
									 x"CC03",x"CC03",x"C403",x"C402",x"C423",x"C423",x"C423",x"C423",x"C423",x"C423",
									 x"C403",x"BC03",x"BC02",x"B402",x"ABC2",x"A342",x"9B01",x"ABE3",x"CDC5",x"F766",
									 x"FFC6",x"FF86",x"FF46",x"FEE5",x"FEC5",x"FEC5",x"FEC6",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE24",x"FE04",x"FDC4",x"FDA4",
									 x"FD83",x"FD43",x"F503",x"FCE2",x"F483",x"EC86",x"E4EB",x"CD72",x"C5D5",x"BDD7",
									 x"C639",x"DEDA",x"EF5D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"EE34",x"F4AA",x"F425",x"EC02",
									 x"F462",x"F483",x"F4C4",x"F504",x"FD24",x"FD44",x"FD64",x"FD84",x"F565",x"FDA7",
									 x"FE6E",x"FF55",x"FF79",x"FF7A",x"FF9A",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF55",
									 x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FEEF",x"FEEE",
									 x"FECE",x"F6AD",x"BCC9",x"59C1",x"5140",x"59A0",x"6A01",x"7241",x"7A61",x"8281",
									 x"82A1",x"8AC1",x"92E2",x"9AE2",x"9B02",x"9B02",x"9B02",x"9B02",x"A322",x"A322",
									 x"A322",x"A322",x"A322",x"9B22",x"9B22",x"9B22",x"9B22",x"92E1",x"92C1",x"8260",
									 x"8260",x"AC45",x"CDE7",x"F74A",x"FF8B",x"FF2A",x"FEC9",x"FE67",x"FE47",x"FE47",
									 x"FE47",x"FE67",x"FE47",x"FE46",x"FE46",x"FE47",x"FE47",x"FE47",x"FE66",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",
									 x"FEA5",x"FEC5",x"EE43",x"BC83",x"8262",x"50C0",x"50E0",x"6160",x"6180",x"6140",
									 x"5940",x"7AC8",x"BD94",x"D6DB",x"E73C",x"E73C",x"E73C",x"E73C",x"EF3D",x"EF3D",
									 x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF7D",x"EF9E",x"FFDF",x"B574",
									 x"41A3",x"3920",x"4980",x"5A00",x"6240",x"7281",x"82C2",x"9301",x"9B21",x"AB42",
									 x"B383",x"BBA2",x"C3C3",x"C3C2",x"C3E2",x"CBE2",x"CC02",x"CC02",x"C402",x"C402",
									 x"C402",x"C422",x"C403",x"C423",x"C423",x"C403",x"BC03",x"BC03",x"B402",x"B3E2",
									 x"ABA2",x"9B42",x"92E1",x"B443",x"DE45",x"F786",x"FFC6",x"FF66",x"FF26",x"FEE5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",
									 x"FE45",x"FE45",x"FE24",x"FE04",x"FDC4",x"FDA4",x"FD84",x"FD23",x"FD03",x"FCC2",
									 x"F483",x"E4A7",x"DD0D",x"CD72",x"C5D6",x"BDF8",x"C659",x"DEDB",x"EF5D",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFDD",x"F696",x"F52D",x"F446",x"EC03",x"F442",x"F463",x"F4C4",x"F504",
									 x"FD04",x"FD24",x"FD44",x"FD64",x"FD65",x"FDA6",x"F62C",x"FF13",x"FF58",x"FF7A",
									 x"FF9A",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",
									 x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FEEF",x"FEEE",x"FEAE",x"E62D",x"9BC7",x"5161",
									 x"4900",x"61C1",x"7241",x"7A61",x"7A81",x"82A1",x"8AC1",x"92C1",x"9B02",x"9B02",
									 x"9B02",x"9B22",x"A322",x"A322",x"A322",x"A342",x"A342",x"A342",x"A342",x"A342",
									 x"A342",x"9B22",x"9B22",x"9301",x"92E1",x"8AA1",x"8281",x"9BA3",x"B4E5",x"EEEA",
									 x"FFAB",x"FF6B",x"FEE9",x"FE88",x"FE47",x"FE47",x"FE67",x"FE67",x"FE47",x"FE46",
									 x"FE46",x"FE47",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FEA5",x"FEC5",x"E604",x"B443",
									 x"7A21",x"50C0",x"58E0",x"6160",x"6180",x"6140",x"5941",x"82C8",x"BD94",x"D6DB",
									 x"E73C",x"E73C",x"E73C",x"E73C",x"EF3D",x"EF3D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",
									 x"EF5D",x"EF5D",x"EF7D",x"EF7D",x"FFBE",x"AD13",x"3942",x"3920",x"49A0",x"5A00",
									 x"6240",x"7281",x"8AC2",x"9301",x"9B21",x"AB42",x"B382",x"BBA2",x"C3C2",x"C3C2",
									 x"C3E2",x"CBE2",x"CC02",x"CC02",x"C402",x"C402",x"C402",x"C422",x"C423",x"C423",
									 x"C403",x"C403",x"BC02",x"BC02",x"B3E3",x"B3C3",x"A382",x"9321",x"9300",x"BCE3",
									 x"EF06",x"FFC6",x"FFA6",x"FF66",x"FF25",x"FEE5",x"FEC5",x"FEC6",x"FEC6",x"FEC5",
									 x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE65",x"FE45",x"FE45",x"FE24",x"FDE4",
									 x"FDC4",x"FDA4",x"FD64",x"FD23",x"FD03",x"FCC3",x"F484",x"E4A8",x"DD2E",x"C573",
									 x"BDD6",x"BE18",x"CE79",x"E6FB",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FEF8",x"F590",
									 x"F467",x"EC03",x"F422",x"F463",x"F4A3",x"F4E4",x"FD04",x"FD24",x"FD44",x"FD64",
									 x"FD65",x"FD85",x"F5E9",x"FED0",x"FF36",x"FF79",x"FF99",x"FF79",x"FF79",x"FF79",
									 x"FF79",x"FF99",x"FF98",x"FF98",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",
									 x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FEEF",x"FEEE",x"F6AD",x"CD4A",x"8304",x"5161",x"5160",x"6201",x"7241",x"7A61",
									 x"8281",x"8AC1",x"8AC1",x"92E1",x"9B02",x"9B22",x"9B22",x"A322",x"A342",x"A342",
									 x"AB42",x"AB42",x"AB42",x"A342",x"AB62",x"A342",x"A342",x"A342",x"9B22",x"9B01",
									 x"9301",x"92C1",x"8A81",x"82A1",x"9382",x"DE89",x"FFCC",x"FF8B",x"FF0A",x"FE88",
									 x"FE67",x"FE47",x"FE47",x"FE67",x"FE47",x"FE46",x"FE46",x"FE47",x"FE47",x"FE47",
									 x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE85",x"FE85",x"FEA5",x"FEC5",x"DDC4",x"AC02",x"7201",x"50E0",x"5900",x"6160",
									 x"6160",x"6140",x"6161",x"82E8",x"BD95",x"D6DB",x"E73C",x"E71C",x"E71C",x"E73C",
									 x"EF3C",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF7D",x"EF5D",
									 x"EF3C",x"9CB0",x"3921",x"3900",x"49A0",x"5A20",x"6A60",x"7281",x"8AE2",x"9301",
									 x"9B21",x"AB62",x"B382",x"BBA2",x"C3C2",x"C3E2",x"C3E2",x"CBE2",x"CC02",x"C402",
									 x"C402",x"C402",x"C402",x"C422",x"C423",x"C403",x"C402",x"BC02",x"BC02",x"B402",
									 x"B3C3",x"ABA3",x"A362",x"9B62",x"9BC1",x"CDC4",x"FF87",x"FFC6",x"FFA6",x"FF45",
									 x"FEE5",x"FEC5",x"FEC6",x"FEC6",x"FEC6",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",
									 x"FE65",x"FE65",x"FE45",x"FE25",x"FE04",x"FDE4",x"FDA4",x"FD84",x"FD63",x"FD03",
									 x"F4E3",x"F4A3",x"EC84",x"DCCA",x"D570",x"C594",x"BDD6",x"C639",x"D69A",x"E71C",
									 x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF5A",x"FDF2",x"F4A9",x"EC24",x"EC22",x"F462",
									 x"F483",x"F4E4",x"FD04",x"FD24",x"FD44",x"FD64",x"FD84",x"FD84",x"FDC8",x"FE8E",
									 x"FEF4",x"FF78",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",x"FF99",x"FF98",x"FF78",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF54",
									 x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"EE6C",x"BCE9",
									 x"7AA3",x"5181",x"5180",x"6A01",x"7261",x"7A61",x"8281",x"8AC1",x"92E1",x"92E1",
									 x"9B02",x"A322",x"A322",x"A342",x"A342",x"A342",x"AB42",x"AB42",x"AB42",x"AB42",
									 x"AB62",x"AB62",x"A362",x"A342",x"A322",x"9B22",x"9B21",x"9B02",x"8AA1",x"7A41",
									 x"82E1",x"DE49",x"FFCC",x"FFAB",x"FF2A",x"FE88",x"FE67",x"FE47",x"FE47",x"FE67",
									 x"FE47",x"FE46",x"FE46",x"FE47",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE86",
									 x"FE86",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FEA5",x"FEC5",x"FEA5",
									 x"DD84",x"A3A2",x"71E0",x"50E0",x"5900",x"6180",x"6160",x"6160",x"6181",x"8B29",
									 x"C5B5",x"D6DB",x"E71C",x"DF1C",x"E71C",x"E73C",x"EF3C",x"EF3D",x"EF5D",x"EF5D",
									 x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5D",x"EF5C",x"DEBA",x"8C0E",x"3921",x"3900",
									 x"51A0",x"6220",x"6A60",x"7A81",x"8AE2",x"9B01",x"9B21",x"AB62",x"B382",x"BBA2",
									 x"C3C2",x"C3E2",x"C3E2",x"CBE2",x"CC02",x"C402",x"C402",x"C402",x"C422",x"C422",
									 x"C422",x"C422",x"C403",x"BC03",x"BC02",x"B3E2",x"B3C3",x"AB82",x"9B21",x"A3E2",
									 x"B4A3",x"DE65",x"FFA7",x"FFC6",x"FF86",x"FF25",x"FEE5",x"FEC5",x"FEC6",x"FEC6",
									 x"FEA6",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE65",x"FE45",x"FE25",
									 x"FE05",x"FDE4",x"FDA4",x"FD84",x"F543",x"FD03",x"F4C2",x"F4A3",x"EC85",x"DCCB",
									 x"CD72",x"BDB5",x"BDD7",x"C659",x"DEBA",x"EF3C",x"FFBF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FF9C",x"FE34",x"F4EB",x"EC25",x"EC22",x"F442",x"F483",x"F4C3",x"FCE3",x"FD04",
									 x"FD44",x"FD64",x"FD84",x"FD84",x"FDC6",x"FE2C",x"FEB2",x"FF58",x"FF99",x"FF9A",
									 x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FEEF",x"FECE",x"EE4C",x"BCC8",x"7281",x"5160",x"5180",x"6A00",
									 x"7261",x"7A61",x"82A1",x"8AC1",x"92E1",x"92E1",x"9B01",x"A322",x"A342",x"A342",
									 x"AB42",x"AB42",x"AB62",x"AB62",x"AB62",x"AB62",x"AB62",x"AB62",x"A342",x"A342",
									 x"A342",x"A321",x"9B21",x"9B02",x"92C2",x"7A01",x"7A60",x"D629",x"FFCD",x"FFAC",
									 x"FF4A",x"FEA8",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE46",x"FE46",x"FE47",
									 x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE85",x"FEA5",x"FEC5",x"F685",x"D544",x"9B82",x"69C0",x"50E0",
									 x"5920",x"6160",x"6160",x"6160",x"69C1",x"936A",x"C5D6",x"D6DB",x"DF1C",x"DF1B",
									 x"E71C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",
									 x"EF5D",x"EF5C",x"CE38",x"7B8C",x"3941",x"3920",x"51C0",x"6220",x"6A60",x"7A81",
									 x"8AE2",x"9B01",x"A341",x"AB62",x"B382",x"BBA2",x"C3C2",x"C3E2",x"C3E2",x"CBE2",
									 x"CC02",x"CC02",x"C402",x"C402",x"C422",x"C422",x"C422",x"C422",x"BC02",x"BC02",
									 x"B402",x"B3E2",x"B3A3",x"AB62",x"9300",x"AC42",x"C564",x"E6E6",x"F7A6",x"FFA6",
									 x"FF46",x"FF06",x"FEC5",x"FEC5",x"FEC6",x"FEC6",x"FEA6",x"FEA5",x"FEA5",x"FEA5",
									 x"FEA5",x"FE85",x"FE65",x"FE45",x"FE45",x"FE05",x"FDE4",x"FDC4",x"FDA4",x"FD64",
									 x"FD43",x"FCE3",x"F4A2",x"F483",x"EC85",x"DD0C",x"CD94",x"BDB6",x"BDF7",x"CE7A",
									 x"DEDB",x"F75C",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"F6B7",x"FD4E",x"EC67",
									 x"EBE2",x"F442",x"F462",x"FCC3",x"F4E3",x"F503",x"FD24",x"FD44",x"FD64",x"FD85",
									 x"FDA6",x"FDE9",x"FE6F",x"FF56",x"FF9A",x"FF9A",x"FF79",x"FF79",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF55",
									 x"FF55",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECF",x"FECF",x"FEAE",
									 x"EE4D",x"BCA8",x"7282",x"51A0",x"5180",x"6A00",x"7241",x"7A61",x"82A1",x"8AC1",
									 x"92E1",x"92E1",x"9B01",x"9B21",x"A342",x"A342",x"AB42",x"AB62",x"AB62",x"AB62",
									 x"AB62",x"AB62",x"AB42",x"AB42",x"A342",x"A342",x"A322",x"9B22",x"9B21",x"9B01",
									 x"92A1",x"7A01",x"7AA1",x"D629",x"FFCC",x"FFAB",x"FF4A",x"FEA8",x"FE67",x"FE67",
									 x"FE47",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE66",x"FE66",x"FE66",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE65",x"FE85",x"FEA5",
									 x"FEC5",x"F665",x"CD04",x"9321",x"69A0",x"50E0",x"6120",x"6160",x"6140",x"6160",
									 x"6A02",x"93AB",x"CDF6",x"D6DB",x"DEFC",x"E71C",x"E71C",x"E73C",x"E73C",x"E73C",
									 x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"EF7D",x"E73C",x"B575",x"6AE9",
									 x"3941",x"4140",x"59C0",x"6241",x"6A60",x"7AA1",x"8AE1",x"9B01",x"A341",x"AB62",
									 x"B382",x"BBA2",x"C3C2",x"C3E2",x"C3E3",x"CC02",x"C402",x"C403",x"C403",x"C403",
									 x"C423",x"C423",x"C423",x"BC03",x"BC02",x"BC02",x"B3E2",x"B3C2",x"A361",x"A342",
									 x"9320",x"C504",x"DE66",x"F786",x"FFA6",x"FF66",x"FF26",x"FF06",x"FEE5",x"FEC5",
									 x"FEC6",x"FEC6",x"FEA6",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE45",x"FE45",
									 x"FE25",x"FE04",x"FDE4",x"FDC4",x"FD84",x"FD44",x"FD24",x"F4E3",x"F4A2",x"F483",
									 x"E487",x"D52E",x"C5D5",x"BDF6",x"BDF7",x"D69A",x"E71C",x"F79D",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFDD",x"F719",x"FDD1",x"ECA9",x"EC03",x"F441",x"F462",x"FCA3",
									 x"F4E3",x"F4E3",x"FD23",x"FD44",x"FD64",x"FD85",x"FD85",x"FDA7",x"FE2C",x"FF15",
									 x"FF79",x"FF7A",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECF",x"FECF",x"FECF",x"F66D",x"C4E9",x"7AC3",x"5180",
									 x"5160",x"6A01",x"7A42",x"7A61",x"82A1",x"8AA1",x"8AE1",x"92E1",x"9B01",x"9B22",
									 x"A342",x"A342",x"A342",x"A342",x"A342",x"A342",x"A342",x"A342",x"AB62",x"A342",
									 x"A342",x"A342",x"A322",x"A302",x"9B01",x"9B00",x"92A1",x"8262",x"8322",x"DE6A",
									 x"FFCD",x"FFAB",x"FF2A",x"FEA7",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FEC5",x"FEE6",x"EE45",x"C4A3",x"8AC0",
									 x"6160",x"5900",x"6140",x"6960",x"6140",x"6180",x"7243",x"93EC",x"CE17",x"D6BA",
									 x"DEFB",x"DEFB",x"E71C",x"E71C",x"E73C",x"E73C",x"E73C",x"E73C",x"E73C",x"E71C",
									 x"E73C",x"E73C",x"EF7D",x"E6FB",x"9CB2",x"5A47",x"4161",x"4960",x"59E0",x"6A41",
									 x"7281",x"7AA0",x"92E1",x"9B02",x"A342",x"AB82",x"B3A2",x"BBA2",x"BBC2",x"C3E2",
									 x"C403",x"C403",x"C403",x"C403",x"C403",x"C403",x"C403",x"C403",x"BC02",x"BC02",
									 x"BBE2",x"BC02",x"B3C2",x"ABA2",x"9B21",x"9B22",x"A3C2",x"D5A6",x"F726",x"FFC6",
									 x"FF87",x"FF46",x"FF06",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA6",
									 x"FEA5",x"FE85",x"FE65",x"FE65",x"FE45",x"FE45",x"FE24",x"FDE4",x"FDE4",x"FDC4",
									 x"FD83",x"FD23",x"FD03",x"F4C3",x"F4A3",x"F4A5",x"E4C9",x"CD50",x"C5D5",x"BE17",
									 x"C618",x"DEDB",x"EF3D",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"F73A",
									 x"FE53",x"ECEB",x"EC04",x"F422",x"F462",x"FCA3",x"F4C3",x"F4E3",x"FD24",x"FD24",
									 x"FD64",x"FD85",x"FD84",x"FDA6",x"F5EA",x"FED2",x"FF58",x"FF7A",x"FF79",x"FF99",
									 x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",
									 x"FF55",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECF",x"F68D",x"CD4A",x"8304",x"5161",x"5161",x"6201",x"7241",x"7A61",
									 x"8281",x"82A1",x"8AC1",x"92E2",x"9302",x"9B22",x"A322",x"A342",x"A342",x"A342",
									 x"A342",x"A342",x"A342",x"A342",x"AB62",x"A342",x"A342",x"A342",x"A322",x"9B02",
									 x"9B01",x"92C1",x"8AA1",x"8AE2",x"93C3",x"DE8A",x"FFCC",x"FF8B",x"FF09",x"FE87",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE66",
									 x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE65",
									 x"FE85",x"FEC5",x"FEE6",x"EE25",x"BC63",x"8260",x"5940",x"5920",x"6140",x"6960",
									 x"5920",x"61A0",x"7284",x"9C2D",x"CE37",x"D6BA",x"DEFB",x"DEFB",x"E71C",x"E71C",
									 x"E71C",x"E71C",x"E71C",x"E71C",x"E71C",x"E71C",x"E71C",x"E73C",x"EF7D",x"E6FB",
									 x"9C70",x"5205",x"4141",x"4960",x"59E0",x"6A41",x"7281",x"82C1",x"9301",x"9B22",
									 x"A342",x"B382",x"BBA2",x"BBC2",x"C3C2",x"C3E2",x"C403",x"C403",x"C403",x"C403",
									 x"C403",x"C403",x"C403",x"BC02",x"BC02",x"BBE2",x"BBE2",x"B3E2",x"B3C2",x"AB82",
									 x"9301",x"9301",x"B444",x"DE46",x"FF86",x"FFC6",x"FF86",x"FF26",x"FEE6",x"FEE5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",
									 x"FE45",x"FE25",x"FE04",x"FDE4",x"FDE4",x"FDC4",x"FD84",x"FD23",x"FCE3",x"F4C3",
									 x"F4A4",x"ECA6",x"DCEB",x"CD71",x"C5D5",x"BE17",x"C638",x"E6DC",x"EF5D",x"F7BE",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",x"F77C",x"FEB7",x"ED4E",x"EC45",x"F423",
									 x"F442",x"FC83",x"F4C3",x"F4E3",x"FD24",x"FD24",x"FD44",x"FD64",x"FD84",x"FDA5",
									 x"FDE8",x"FE8F",x"FF56",x"FF7A",x"FF9A",x"FF99",x"FF79",x"FF79",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF35",x"FF35",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FEAE",x"E5EB",
									 x"9BC6",x"5161",x"4920",x"61C0",x"7241",x"7A41",x"8281",x"82A1",x"8AC2",x"92E2",
									 x"92E2",x"9B02",x"9B22",x"A342",x"A322",x"A322",x"A322",x"A342",x"A342",x"A342",
									 x"A342",x"A342",x"A322",x"A322",x"9B21",x"9B02",x"9AE2",x"8AA1",x"8260",x"9383",
									 x"ACA5",x"E6CA",x"FFAC",x"FF6B",x"FEE9",x"FE87",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FE84",x"FEC4",x"FEE6",x"E605",
									 x"AC03",x"7A21",x"5900",x"5920",x"6160",x"6960",x"6140",x"61A1",x"7AE6",x"A48F",
									 x"CE58",x"D6BA",x"DEFB",x"DEFB",x"E71C",x"E71C",x"E71C",x"E71C",x"E71C",x"E71C",
									 x"E71C",x"E71C",x"E71C",x"E73C",x"EF9E",x"DEDA",x"8C2F",x"41A3",x"4160",x"51A0",
									 x"59E0",x"6A41",x"7281",x"82C1",x"9301",x"A322",x"AB42",x"B383",x"BBA2",x"BBC2",
									 x"C3C2",x"C3E2",x"C3E2",x"C403",x"C403",x"C3E2",x"C402",x"C402",x"C403",x"BC02",
									 x"BBE2",x"BBE2",x"B3C2",x"B3C2",x"B3C3",x"A362",x"8B00",x"9361",x"C525",x"EEE6",
									 x"FFC6",x"FFA6",x"FF46",x"FF06",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE24",x"FE04",x"FDC4",
									 x"FDC4",x"FDA4",x"FD64",x"FD23",x"FCE3",x"F4A3",x"EC84",x"E4A8",x"D50E",x"C573",
									 x"BDD6",x"C637",x"CE79",x"E71C",x"F77E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"F7BE",x"FF5A",x"EDD1",x"E467",x"EC23",x"F422",x"FC62",x"F4A3",x"FCE4",
									 x"FD04",x"FD24",x"FD44",x"FD64",x"FD85",x"FD85",x"FDA6",x"FE4C",x"FF14",x"FF79",
									 x"FF9A",x"FF79",x"FF79",x"FF79",x"FF79",x"FF79",x"FF78",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF55",x"FF55",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECF",x"FEEF",x"FEEE",x"FECE",x"F6AE",x"BCC9",x"6A02",x"5160",x"59C0",
									 x"6A21",x"7221",x"7A61",x"8281",x"82A1",x"8AC1",x"8AC1",x"92E1",x"9B02",x"9B02",
									 x"9B02",x"9B02",x"A322",x"A322",x"A322",x"A322",x"A322",x"9B22",x"9B22",x"9B22",
									 x"9B01",x"9AE1",x"92C2",x"8261",x"7A80",x"B4A5",x"D608",x"F74A",x"FF8B",x"FF2A",
									 x"FEC8",x"FE67",x"FE47",x"FE47",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE85",x"FE85",x"FE84",x"FEC4",x"FEE6",x"E5C4",x"A382",x"69C1",x"50C0",x"5940",
									 x"6960",x"6940",x"5920",x"61C2",x"8349",x"ACF2",x"D679",x"D6BA",x"DEDB",x"DEDB",
									 x"DEFB",x"E71C",x"E71C",x"E71C",x"DEFB",x"E71C",x"E71C",x"E71C",x"E71C",x"E73C",
									 x"EF5D",x"D699",x"7B8C",x"3941",x"4180",x"51A0",x"6200",x"7261",x"7A81",x"82E1",
									 x"9B21",x"A322",x"AB42",x"B382",x"BBA2",x"C3C2",x"C3C2",x"C3E2",x"C3E2",x"C403",
									 x"C403",x"C3E2",x"C402",x"C402",x"C402",x"BBE2",x"BBE2",x"BBC2",x"B3C2",x"ABA2",
									 x"A362",x"9B21",x"9BA1",x"AC42",x"DE47",x"FF87",x"FFC6",x"FF86",x"FF26",x"FEE5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE65",x"FE45",x"FE24",x"FE04",x"FDE4",x"FDC4",x"FDA4",x"FDA4",x"FD44",x"FD03",
									 x"FCC3",x"F483",x"EC85",x"DCCB",x"D551",x"C5B4",x"BDD6",x"C658",x"D6BA",x"EF3D",
									 x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"F634",
									 x"ECC9",x"F444",x"F422",x"FC42",x"F483",x"F4C3",x"F4E4",x"FD04",x"FD24",x"FD44",
									 x"FD65",x"FD64",x"FD85",x"FE0A",x"FEF2",x"FF57",x"FF79",x"FF79",x"FF79",x"FF79",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF57",
									 x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF35",
									 x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FEEE",
									 x"FEEE",x"FEEE",x"D58B",x"9345",x"7262",x"59A0",x"59C1",x"6A00",x"7220",x"7A61",
									 x"8281",x"8AA1",x"8AC1",x"92C1",x"92E1",x"92E1",x"9B02",x"9B02",x"9B02",x"9B02",
									 x"9B02",x"9B02",x"9B22",x"9B01",x"9B02",x"9302",x"92E1",x"92C1",x"8A61",x"7A40",
									 x"8B21",x"CDA8",x"EF0A",x"FF8A",x"FF4A",x"FEE9",x"FEA8",x"FE67",x"FE47",x"FE47",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE66",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE66",x"FE85",x"FEA4",x"FEC4",
									 x"FEE6",x"DDA4",x"9B42",x"6161",x"48A0",x"6140",x"6980",x"6961",x"5900",x"61C3",
									 x"838B",x"AD34",x"D67A",x"D6BB",x"DEDB",x"DEDB",x"DEFB",x"DEFB",x"DEFB",x"DEFB",
									 x"DEFB",x"DEFB",x"E71C",x"E71C",x"E71C",x"E73C",x"E73C",x"CE58",x"732A",x"3100",
									 x"4980",x"51C0",x"6201",x"7262",x"7AA1",x"8AE1",x"9B22",x"A322",x"AB42",x"B382",
									 x"BBA2",x"C3C2",x"C3C2",x"C3E2",x"C3E2",x"C3E2",x"C3E2",x"C3E2",x"C3E2",x"C3E2",
									 x"BBE2",x"BBE2",x"BBC2",x"B3C2",x"B3A2",x"AB82",x"9B01",x"9321",x"AC62",x"C563",
									 x"EF07",x"FFC7",x"FFA5",x"FF45",x"FF05",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE24",x"FE04",
									 x"FDE4",x"FDC3",x"FDA4",x"FD84",x"F524",x"F4E3",x"F4C2",x"F482",x"EC86",x"DCED",
									 x"D593",x"C5D6",x"BDF7",x"CE79",x"DEDB",x"EF5E",x"FFBF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"F696",x"F52D",x"F466",x"F423",x"F442",
									 x"F483",x"F4A4",x"F4E4",x"F504",x"FD24",x"FD44",x"FD64",x"FD84",x"FD84",x"FDE8",
									 x"FEAF",x"FF35",x"FF58",x"FF79",x"FF79",x"FF79",x"FF78",x"FF79",x"FF78",x"FF78",
									 x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FF12",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FEEE",x"EE2C",x"BCA8",
									 x"9344",x"59A0",x"5981",x"69E1",x"7221",x"7A61",x"7A61",x"8281",x"8AA1",x"8AC1",
									 x"92C1",x"92E1",x"9301",x"9B01",x"9B02",x"9AE2",x"9B02",x"9B02",x"9B02",x"9AE2",
									 x"9AE2",x"92E2",x"92A1",x"8A61",x"7A00",x"82A1",x"AC64",x"DE89",x"FF8B",x"FF8A",
									 x"FF29",x"FEC8",x"FE87",x"FE47",x"FE47",x"FE47",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FEC4",x"FEC6",x"D544",x"9302",x"6141",
									 x"4880",x"6140",x"6980",x"6960",x"5900",x"61C3",x"8BAC",x"B555",x"D69B",x"DEDB",
									 x"D6BB",x"DEDB",x"DEFB",x"DEFB",x"DEFB",x"DEFB",x"E71C",x"DEFC",x"E71C",x"E71C",
									 x"E71B",x"E73C",x"DF1B",x"C5F6",x"6B09",x"3100",x"4980",x"51C0",x"6221",x"7281",
									 x"7AA1",x"8AE1",x"9B22",x"A322",x"AB62",x"B382",x"BBA2",x"C3C2",x"C3C2",x"C3E2",
									 x"C3E2",x"C3E2",x"C3E2",x"C3E2",x"C3E2",x"C3E2",x"BBE2",x"BBE2",x"B3C2",x"B3C2",
									 x"AB82",x"A362",x"9B01",x"9B41",x"C523",x"DE65",x"F787",x"FFC7",x"FF86",x"FF25",
									 x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",
									 x"FE85",x"FE65",x"FE45",x"FE45",x"FE24",x"FE05",x"FDE4",x"FDA4",x"FD84",x"F564",
									 x"F523",x"F4E3",x"F4A2",x"F463",x"E4A8",x"DD2F",x"CD73",x"C5D6",x"BE18",x"CE99",
									 x"DEFB",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FF19",x"F5B0",x"F489",x"F404",x"F402",x"F463",x"F4A4",x"F4C4",x"F504",
									 x"FD24",x"F544",x"FD64",x"FD84",x"F584",x"FDA6",x"FE4C",x"FED3",x"FF57",x"FF99",
									 x"FF9A",x"FF79",x"FF58",x"FF59",x"FF79",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",
									 x"FF77",x"FF77",x"FF57",x"FF57",x"FF56",x"FF56",x"FF36",x"FF36",x"FF36",x"FF55",
									 x"FF55",x"FF35",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FF11",
									 x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FEEF",x"FECE",x"FECE",x"FEEE",x"FECD",x"E60B",x"BCE8",x"82C3",x"61C0",x"5980",
									 x"61C0",x"7201",x"7A61",x"7A61",x"8281",x"8AA2",x"8AC1",x"8AC1",x"92C1",x"92E1",
									 x"92E2",x"92E2",x"92E2",x"92E2",x"92C1",x"92C2",x"92A2",x"8AA1",x"8261",x"8242",
									 x"82A2",x"9BC3",x"D608",x"F74B",x"FF8A",x"FF49",x"FEC8",x"FE88",x"FE47",x"FE27",
									 x"FE47",x"FE47",x"FE67",x"FE47",x"FE47",x"FE46",x"FE47",x"FE47",x"FE46",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",
									 x"FE86",x"FEA4",x"FEA5",x"CCE4",x"8AC1",x"5920",x"4880",x"6141",x"6980",x"6960",
									 x"5900",x"69E4",x"93CD",x"BD95",x"D6BA",x"D6BA",x"D6BA",x"D6BA",x"DEDB",x"DEFB",
									 x"DEFB",x"DEFB",x"DEFC",x"DEFC",x"E71C",x"E71C",x"E71B",x"E73C",x"CE78",x"A513",
									 x"62A8",x"3900",x"4980",x"59C0",x"6241",x"7281",x"82A1",x"92C1",x"A301",x"AB42",
									 x"AB62",x"B382",x"BBA2",x"BBC2",x"C3C2",x"C3C2",x"C3E2",x"C3E2",x"C3E2",x"C3E2",
									 x"C3E2",x"BBE3",x"BBC3",x"B3C3",x"B3E2",x"ABA2",x"A363",x"9B21",x"9321",x"AC22",
									 x"D605",x"EF06",x"FF87",x"FF86",x"FF45",x"FF05",x"FEE5",x"FEE5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",x"FE25",
									 x"FE05",x"FE05",x"FDE4",x"FDA4",x"FD84",x"FD43",x"F503",x"F4C3",x"F4A3",x"F484",
									 x"E4EA",x"D551",x"CD94",x"C5F7",x"BE59",x"D6BA",x"E73C",x"F7DF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF7B",x"FE34",x"F4EB",
									 x"F425",x"F402",x"F462",x"F483",x"F4C3",x"F4E4",x"F524",x"F524",x"FD44",x"FD85",
									 x"FD85",x"FDA5",x"FDE9",x"FE6F",x"FF15",x"FF79",x"FF9A",x"FF79",x"FF58",x"FF59",
									 x"FF78",x"FF78",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",
									 x"FF56",x"FF56",x"FF36",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF55",x"FF54",
									 x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FF11",x"FEF0",x"FEF0",x"FED0",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",
									 x"FEEE",x"F6AE",x"EE2C",x"BCC9",x"8B03",x"6A00",x"61C0",x"61C1",x"7223",x"7222",
									 x"7A42",x"8261",x"8281",x"82A1",x"8AA1",x"8AA1",x"8AA2",x"8AC2",x"8AC1",x"8AC1",
									 x"8AA1",x"8A81",x"8A62",x"8262",x"7240",x"8B02",x"B485",x"CD87",x"F70B",x"FF6B",
									 x"FF49",x"FEE9",x"FEA8",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE46",x"FE47",x"FE47",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE86",x"FEA5",x"FE85",x"C4A4",
									 x"8281",x"5920",x"50A0",x"6140",x"6980",x"6160",x"5900",x"6A05",x"9BEE",x"BDB6",
									 x"D6BA",x"D69A",x"D69A",x"D6BA",x"DEDB",x"DEDB",x"DEDB",x"DEFB",x"DEFB",x"DEFB",
									 x"DEFB",x"DEFB",x"E71C",x"E73C",x"BDB6",x"8C0E",x"5226",x"3920",x"51A0",x"59E0",
									 x"6A41",x"7A81",x"82A1",x"92E1",x"A322",x"AB42",x"AB42",x"B382",x"BBA2",x"BBC2",
									 x"C3C2",x"C3C2",x"C3E2",x"C3E2",x"C3E2",x"BBE2",x"BBE2",x"BBE2",x"B3C2",x"B3C2",
									 x"B3C2",x"AB82",x"9B22",x"9301",x"9BA1",x"C564",x"EF07",x"FFA7",x"FFA7",x"FF66",
									 x"FF25",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",
									 x"FE65",x"FE65",x"FE65",x"FE44",x"FE24",x"FE24",x"FE04",x"FDE4",x"FDC4",x"FD83",
									 x"FD63",x"F523",x"F503",x"F4C3",x"EC83",x"EC86",x"DD0C",x"CD92",x"BDB5",x"BDF7",
									 x"CE7A",x"DEFB",x"EF7D",x"F7DF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"FEB7",x"F56F",x"EC67",x"F402",x"F442",x"F483",
									 x"F4A3",x"F4C4",x"F504",x"F524",x"FD44",x"FD65",x"FD85",x"FD85",x"FDA7",x"FE0B",
									 x"FED2",x"FF78",x"FF7A",x"FF7A",x"FF58",x"FF58",x"FF58",x"FF78",x"FF78",x"FF78",
									 x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF55",x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",
									 x"FEF1",x"FF11",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FEEF",x"FECE",x"FECE",x"FECE",x"FECD",x"FECE",x"FEAD",x"E60B",
									 x"BCC7",x"9BC5",x"7AC2",x"61E1",x"61A1",x"61E1",x"6A01",x"7241",x"7A61",x"8281",
									 x"8281",x"8281",x"8281",x"8281",x"8281",x"8261",x"7A61",x"7A21",x"7A41",x"7A82",
									 x"8B63",x"BD06",x"DE28",x"EEC9",x"FF2A",x"FF29",x"FEC8",x"FE88",x"FE67",x"FE67",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE47",x"FE47",
									 x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE85",x"FEA6",x"FEA5",x"F645",x"BC43",x"7A41",x"5920",x"50C0",x"6160",
									 x"6980",x"6140",x"5920",x"6A05",x"9C0E",x"BDD6",x"D6DA",x"CEBA",x"D69A",x"D6BA",
									 x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"DEFB",x"DEDB",x"DEFB",x"DEFB",x"E73C",x"EF5D",
									 x"B554",x"734B",x"51E4",x"4140",x"51A0",x"6200",x"6A41",x"7AA2",x"8AC1",x"9AE1",
									 x"A322",x"AB42",x"B362",x"BB82",x"BBA2",x"C3C2",x"C3C2",x"C3E2",x"C3E2",x"C3E2",
									 x"BBE2",x"BBC2",x"BBC2",x"BBC2",x"B3C2",x"ABA2",x"AB82",x"A342",x"9B22",x"9B41",
									 x"AC41",x"D645",x"F766",x"FFA7",x"FF66",x"FF26",x"FF05",x"FEE5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE44",
									 x"FE24",x"FE04",x"FDE4",x"FDC4",x"FDA4",x"FD63",x"FD42",x"F522",x"F4E3",x"F4A3",
									 x"ECA4",x"E4A9",x"D54F",x"C5D4",x"B5D6",x"C618",x"D69A",x"E73C",x"F79D",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FF5B",x"F5F3",x"F4CA",x"F403",x"F422",x"F463",x"F4A3",x"F4C3",x"F4E4",x"F504",
									 x"FD44",x"FD65",x"FD65",x"FD85",x"FD86",x"FDC9",x"FE90",x"FF56",x"FF79",x"FF79",
									 x"FF79",x"FF58",x"FF58",x"FF58",x"FF78",x"FF78",x"FF77",x"FF77",x"FF77",x"FF77",
									 x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF55",
									 x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FF11",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FEEF",x"FECE",
									 x"FECE",x"FECE",x"FEAD",x"FECD",x"FEED",x"FECD",x"EE4B",x"DDAA",x"AC66",x"82E2",
									 x"6A21",x"6A21",x"6A20",x"7220",x"7220",x"7220",x"7241",x"7A41",x"7A61",x"7A41",
									 x"7A41",x"7A61",x"7A61",x"7A81",x"82E2",x"9362",x"BD06",x"E669",x"FF2A",x"FF4A",
									 x"FF09",x"FEA8",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE46",x"FE47",x"FE47",x"FE46",x"FE66",x"FE66",x"FE66",
									 x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FEA6",x"F684",
									 x"EE04",x"B403",x"7201",x"5921",x"5900",x"6160",x"6960",x"6140",x"5940",x"7245",
									 x"9C2E",x"C5D6",x"D6BA",x"CE9A",x"D69A",x"DEBB",x"DEDB",x"DEDB",x"DEDB",x"DEDB",
									 x"DEFB",x"DEDB",x"DEFB",x"DEFB",x"E71C",x"EF5D",x"A4F2",x"62A8",x"49A3",x"4960",
									 x"59C0",x"6220",x"7241",x"82A2",x"8AC1",x"9AE1",x"AB22",x"AB42",x"B362",x"BB82",
									 x"BBA2",x"C3C2",x"C3E2",x"C3E2",x"C3E2",x"BBE2",x"BBC2",x"BBC2",x"BBC2",x"B3C2",
									 x"B3A2",x"B3A2",x"A362",x"9B22",x"9321",x"A3C1",x"BD23",x"EF26",x"FFA6",x"FFA6",
									 x"FF46",x"FF06",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE65",x"FE45",x"FE24",x"FE04",x"FE04",x"FDE4",x"FDC4",
									 x"FDA4",x"FD63",x"FD23",x"FD02",x"F4C3",x"ECA4",x"ECA6",x"DCCB",x"CD71",x"BDF6",
									 x"B5F7",x"C638",x"DEDB",x"EF5C",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF9D",x"FE97",x"FD6D",x"F425",
									 x"F422",x"F443",x"F463",x"F4A3",x"F4E3",x"FD04",x"FD24",x"FD44",x"FD85",x"FD85",
									 x"FD85",x"F5C8",x"F62C",x"FEF3",x"FF77",x"FF79",x"FF79",x"FF78",x"FF58",x"FF58",
									 x"FF58",x"FF77",x"FF77",x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",x"FF56",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",
									 x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FF12",x"FEF1",x"FEF1",x"FF11",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FECD",
									 x"FECD",x"FECD",x"FECD",x"F6AD",x"EE4C",x"D58A",x"BCC8",x"AC26",x"9384",x"82E3",
									 x"7A82",x"7241",x"6A00",x"69E0",x"6A00",x"7240",x"82C2",x"9343",x"AC05",x"BCE6",
									 x"D5A8",x"E628",x"F6C9",x"FF29",x"FF28",x"FEE8",x"FEA8",x"FE68",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",
									 x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE85",x"FEA6",x"F684",x"E5C4",x"A362",x"69A0",x"5900",
									 x"5901",x"6160",x"6960",x"6140",x"69A1",x"7AA6",x"A46F",x"C5F7",x"D69A",x"CE9A",
									 x"D69A",x"D6BA",x"DEDB",x"DEDB",x"DEDB",x"DEDB",x"DEDA",x"DEDA",x"DEDB",x"DEDB",
									 x"E71C",x"E73D",x"9470",x"49E5",x"4161",x"4980",x"59E0",x"6220",x"7261",x"82A2",
									 x"92C1",x"9B01",x"AB42",x"AB42",x"B362",x"BB82",x"BBA2",x"BBC2",x"C3C2",x"C3E2",
									 x"BBE2",x"BBC2",x"BBC2",x"BBC2",x"B3C2",x"B3A2",x"B382",x"B362",x"A321",x"9301",
									 x"9B82",x"BCE4",x"DE66",x"FFA8",x"FF86",x"FF66",x"FF06",x"FEE5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEC6",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE45",
									 x"FE45",x"FE24",x"FE04",x"FE04",x"FDE4",x"FDA4",x"FDA4",x"F544",x"FD23",x"FCE3",
									 x"F4A3",x"EC85",x"ECA7",x"D50D",x"CD92",x"C5F7",x"BE18",x"CE79",x"E71C",x"F77D",
									 x"FFDE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFBE",x"FF1A",x"FDF1",x"EC66",x"F424",x"F423",x"F443",x"F483",
									 x"F4E4",x"FCE3",x"FD24",x"FD44",x"FD65",x"FD84",x"F585",x"F5A6",x"F5E9",x"FEB0",
									 x"FF56",x"FF79",x"FF79",x"FF78",x"FF58",x"FF58",x"FF58",x"FF57",x"FF77",x"FF77",
									 x"FF77",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF56",x"FF55",
									 x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FF11",
									 x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FECC",x"FECC",x"FECD",
									 x"FECD",x"FEAC",x"EE4B",x"DDAA",x"C508",x"BCA7",x"B446",x"AC06",x"A3C5",x"9BA4",
									 x"A3A3",x"AC04",x"B465",x"C4E6",x"D567",x"E628",x"FECA",x"FEE9",x"FF09",x"FF08",
									 x"FEC8",x"FEA8",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",
									 x"FEC6",x"F665",x"DD64",x"9AE1",x"5940",x"5900",x"6120",x"6160",x"6960",x"6140",
									 x"69C1",x"7AE6",x"A4AF",x"C5F7",x"CE9A",x"CE7B",x"D69A",x"D6BA",x"D6BA",x"DEDB",
									 x"DEDB",x"DEDB",x"DEDA",x"DEDA",x"DEFB",x"D6DB",x"E71C",x"E71C",x"8C0E",x"4183",
									 x"4140",x"4980",x"6200",x"6A40",x"7A81",x"8AC2",x"92C2",x"A301",x"AB42",x"AB62",
									 x"B362",x"BB82",x"BBA2",x"BBA2",x"BBC2",x"BBC2",x"BBC2",x"BBC2",x"BBC2",x"B3A2",
									 x"B3A2",x"B382",x"AB62",x"A342",x"9B01",x"9B62",x"B463",x"D5E5",x"F727",x"FFA7",
									 x"FF66",x"FF45",x"FF05",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC6",x"FEA5",
									 x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE25",x"FE24",x"FE04",x"FDE4",
									 x"FDC4",x"FDA4",x"FD84",x"FD44",x"FD03",x"FCC3",x"F483",x"EC85",x"E4EA",x"CD50",
									 x"C594",x"C5F7",x"C618",x"D69A",x"E75C",x"F79D",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",x"FF9C",
									 x"FE75",x"ECA9",x"EC25",x"F403",x"F423",x"F483",x"F4C4",x"FCE3",x"FD04",x"FD24",
									 x"FD44",x"FD64",x"FD84",x"FDA5",x"F5C7",x"FE6C",x"FF14",x"FF59",x"FF7A",x"FF79",
									 x"FF58",x"FF58",x"FF58",x"FF57",x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF54",
									 x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FF11",x"FEF0",x"FEF0",x"FED0",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FECC",x"FECD",x"FEAC",x"FEAD",x"FEAC",x"F68C",x"F66B",
									 x"EE4B",x"EE4B",x"EE2B",x"EE2B",x"EE2A",x"EE2A",x"EE09",x"EE08",x"EE28",x"F648",
									 x"F668",x"FEA8",x"FEA9",x"FEA9",x"FEC8",x"FE88",x"FE87",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",
									 x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FEC6",x"EE45",x"D505",x"9280",
									 x"5100",x"5900",x"6140",x"6961",x"6161",x"6141",x"6A02",x"8328",x"A4D0",x"C617",
									 x"CE9A",x"D67B",x"D69A",x"D6BA",x"D6BA",x"D6BA",x"D6BA",x"DEDB",x"D6BA",x"D6DA",
									 x"D6DB",x"D6FB",x"DEFB",x"D679",x"7B8C",x"3962",x"4140",x"51A0",x"6201",x"6A41",
									 x"7A81",x"8AC2",x"92E2",x"A302",x"AB42",x"AB62",x"B362",x"BB82",x"BBA2",x"BBA2",
									 x"BBC2",x"BBC2",x"BBC2",x"BBC2",x"B3A2",x"B3A2",x"B382",x"AB62",x"AB43",x"9B22",
									 x"9301",x"A3E2",x"C564",x"E6E5",x"FFA7",x"FFA7",x"FF46",x"FF26",x"FF05",x"FEC5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA6",x"FEA6",x"FE85",x"FE85",x"FE65",x"FE45",
									 x"FE45",x"FE45",x"FE25",x"FE05",x"FDE4",x"FDC4",x"FDC4",x"FDA4",x"FD64",x"FD23",
									 x"FD03",x"FCC2",x"F483",x"E487",x"DD2D",x"C5B3",x"C5B5",x"BDF7",x"C679",x"DEDB",
									 x"EF7E",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FF19",x"F54E",x"F487",x"F424",
									 x"F422",x"F442",x"F4A3",x"FCC3",x"FCE4",x"FD24",x"FD44",x"FD44",x"FD85",x"FD85",
									 x"FDA5",x"FE0A",x"FEB0",x"FF16",x"FF79",x"FF79",x"FF78",x"FF58",x"FF58",x"FF57",
									 x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",
									 x"FEF1",x"FF11",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FECC",x"FECC",x"FECB",x"FECB",x"FECB",
									 x"FECB",x"FECA",x"FEA9",x"FEA9",x"FEA8",x"FEA7",x"FEA7",x"FEA8",x"FE88",x"FE88",
									 x"FE88",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE85",x"FEC6",x"EE05",x"C484",x"8220",x"48A0",x"58E0",x"6961",x"6961",
									 x"6140",x"6140",x"7243",x"8BAA",x"AD32",x"C637",x"CE7A",x"D69A",x"D69A",x"D69A",
									 x"D6BA",x"D6BA",x"D6BA",x"D6BA",x"D6BA",x"D6BA",x"DEDB",x"DEDB",x"D69A",x"B555",
									 x"6AC8",x"3941",x"4160",x"59C0",x"6200",x"6A61",x"7A81",x"8AC2",x"92E2",x"A302",
									 x"AB42",x"AB62",x"B382",x"BBA2",x"BBA2",x"BBA2",x"BBC2",x"BBC2",x"BBC2",x"B3A2",
									 x"B3A2",x"B382",x"AB62",x"A342",x"9AE2",x"9B02",x"9BA1",x"C564",x"EEC6",x"F767",
									 x"FFC7",x"FF66",x"FF26",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",
									 x"FEA5",x"FEA5",x"FE85",x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE25",x"FE04",
									 x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD63",x"FD03",x"FCE3",x"FCA3",x"F484",x"E4C9",
									 x"D56F",x"C5D5",x"C5D7",x"C619",x"D69A",x"E71C",x"F79E",x"FFDF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"F7FF",x"FFFF",x"FF7C",x"F613",x"F50A",x"EC25",x"F402",x"F422",x"F463",x"F4A3",
									 x"FCE3",x"FD04",x"FD24",x"FD44",x"FD65",x"FD85",x"FD85",x"FDE7",x"FE4C",x"FED2",
									 x"FF57",x"FF79",x"FF58",x"FF58",x"FF58",x"FF57",x"FF77",x"FF77",x"FF77",x"FF57",
									 x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF36",x"FF56",x"FF55",x"FF55",x"FF55",
									 x"FF55",x"FF54",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FF12",x"FF12",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FECC",x"FEAC",x"FEAB",x"FEAB",x"FEAB",
									 x"FE8B",x"FEAB",x"FEAB",x"FEAB",x"FEAB",x"FEAB",x"FEAA",x"FE89",x"FE89",x"FE67",
									 x"FE67",x"FE46",x"FE46",x"FE67",x"FE68",x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FE65",x"FEA5",x"FEC6",x"E5C5",
									 x"BC24",x"71A0",x"4880",x"58E0",x"6961",x"6960",x"6140",x"6160",x"72A6",x"9C2D",
									 x"BD94",x"C638",x"CE7A",x"D69A",x"D69A",x"D69A",x"D6BA",x"D6BA",x"D6BA",x"D6BA",
									 x"D69A",x"D6BA",x"DEDC",x"E6FC",x"CE38",x"8C2F",x"5225",x"3940",x"4980",x"59E0",
									 x"6220",x"6A61",x"7A81",x"8AE2",x"92E2",x"A322",x"AB42",x"B362",x"B382",x"BBA2",
									 x"BBA2",x"BBA2",x"BBC2",x"BBC2",x"BBC2",x"B3A2",x"B382",x"AB62",x"A342",x"A322",
									 x"92E1",x"9B82",x"B481",x"E665",x"F786",x"FFA6",x"FF86",x"FF25",x"FF05",x"FEE5",
									 x"FEC5",x"FEC5",x"FEA5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE65",
									 x"FE65",x"FE45",x"FE25",x"FE25",x"FE05",x"FDE5",x"FDC4",x"FDC4",x"FD84",x"FD64",
									 x"FD43",x"FCE3",x"F4C3",x"F484",x"EC86",x"DD0D",x"CD92",x"BDD6",x"C5F8",x"CE5A",
									 x"DEDB",x"EF5C",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FEB7",
									 x"F58E",x"E467",x"EC03",x"FC22",x"F463",x"F4A3",x"FCE3",x"FD03",x"FD24",x"FD24",
									 x"FD45",x"FD65",x"FD85",x"FDC6",x"FE09",x"FE6E",x"FF34",x"FF78",x"FF58",x"FF58",
									 x"FF58",x"FF78",x"FF77",x"FF77",x"FF77",x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF56",x"FF55",x"FF55",x"FF55",x"FF55",x"FF54",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAB",x"FE8B",x"FEAB",
									 x"FEAB",x"FE8B",x"FE8B",x"FE8A",x"FE69",x"FE68",x"FE47",x"FE47",x"FE67",x"FE68",
									 x"FE48",x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",x"FE66",x"FE65",
									 x"FE65",x"FE65",x"FE85",x"FEA5",x"FEA6",x"DDA5",x"B404",x"71A1",x"4880",x"5900",
									 x"6961",x"6960",x"5920",x"5941",x"7AE8",x"A490",x"BDB6",x"CE5A",x"CE7A",x"D679",
									 x"D679",x"D69A",x"D69A",x"D6BA",x"D6BA",x"D6BA",x"D6BA",x"D69A",x"DEDC",x"E6FC",
									 x"CE17",x"7B8C",x"49E3",x"4160",x"4980",x"59E0",x"6220",x"7261",x"8281",x"92E2",
									 x"9AE1",x"A322",x"AB42",x"B361",x"BB82",x"BBA2",x"BBA2",x"BBA2",x"BBA2",x"BBA2",
									 x"B3A2",x"B382",x"AB62",x"A342",x"9B22",x"9B01",x"9341",x"B463",x"CDA4",x"F746",
									 x"FFC6",x"FFA6",x"FF46",x"FF05",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",
									 x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE25",x"FE25",
									 x"FE05",x"FDE5",x"FDC4",x"FDA4",x"FD84",x"FD64",x"FD23",x"FCC3",x"F4A4",x"EC85",
									 x"E488",x"D550",x"C5B5",x"BDD6",x"C618",x"D69A",x"DEFB",x"F77D",x"FFDF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FF5A",x"F632",x"E4CA",x"F424",x"FC03",
									 x"F443",x"F4A3",x"F4E3",x"F503",x"F504",x"FD25",x"FD65",x"FD85",x"FD85",x"FDA5",
									 x"FDC7",x"FE2B",x"FEB0",x"FF36",x"FF58",x"FF78",x"FF78",x"FF57",x"FF57",x"FF57",
									 x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF35",
									 x"FF35",x"FF55",x"FF35",x"FF54",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8B",x"FE8A",
									 x"FE69",x"FE68",x"FE47",x"FE47",x"FE67",x"FE47",x"FE47",x"FE48",x"FE47",x"FE47",
									 x"FE47",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE66",x"FE66",x"FE65",x"FE45",x"FE65",x"FE85",x"FEA5",
									 x"F665",x"D564",x"A363",x"6141",x"50A0",x"5900",x"6980",x"6960",x"5920",x"5941",
									 x"832A",x"A4D2",x"BDF8",x"CE7A",x"CE59",x"CE58",x"CE79",x"D69A",x"D69A",x"D69A",
									 x"D69A",x"D69A",x"D6BA",x"CE9A",x"D6DC",x"E71C",x"BDD6",x"62C8",x"3961",x"4180",
									 x"4980",x"6200",x"6A41",x"7281",x"82A1",x"92E2",x"9AE1",x"A321",x"B341",x"B361",
									 x"B382",x"BB82",x"BB82",x"BB82",x"B382",x"B382",x"B381",x"AB61",x"A342",x"A322",
									 x"92E1",x"9301",x"AC03",x"CD85",x"EEC6",x"FF87",x"FFA6",x"FF26",x"FF06",x"FEE5",
									 x"FEC5",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",
									 x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE05",x"FDE4",x"FDE5",x"FDC4",x"FDA4",
									 x"FD64",x"FD23",x"FCE3",x"FCA3",x"F484",x"EC86",x"E4CA",x"D592",x"C5D7",x"BDD6",
									 x"CE39",x"DEDB",x"EF5C",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFBD",x"FED7",x"F5AF",x"F467",x"F402",x"F422",x"F483",x"F4C3",x"F4E3",
									 x"F504",x"F524",x"F545",x"F565",x"F565",x"FD85",x"FDA5",x"FDE8",x"FE6E",x"FEF4",
									 x"FF57",x"FF78",x"FF58",x"FF58",x"FF57",x"FF57",x"FF57",x"FF57",x"FF57",x"FF56",
									 x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF35",x"FF35",x"FF35",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE89",x"FE69",x"FE68",x"FE67",x"FE66",
									 x"FE66",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",
									 x"FE66",x"FE65",x"FE45",x"FE65",x"FEA5",x"FEA5",x"F645",x"CCE3",x"9302",x"6141",
									 x"50A0",x"6100",x"6960",x"6160",x"5940",x"5962",x"836A",x"ACF3",x"BDF8",x"CE5A",
									 x"CE39",x"CE58",x"CE79",x"CE79",x"D69A",x"D69A",x"D69A",x"D69A",x"D699",x"D6BA",
									 x"D6DC",x"DEDB",x"B553",x"5245",x"3120",x"4180",x"51A0",x"6220",x"7261",x"7281",
									 x"82A1",x"92E2",x"9B01",x"A321",x"B341",x"B361",x"B382",x"B382",x"B382",x"B382",
									 x"B382",x"B381",x"AB41",x"A342",x"A322",x"9B02",x"9301",x"9BA2",x"CD85",x"EEC7",
									 x"FF88",x"FFA7",x"FF45",x"FF05",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",
									 x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE24",
									 x"FE25",x"FE04",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD44",x"FD23",x"FCC3",x"F4A3",
									 x"F484",x"ECA7",x"E50E",x"CD94",x"BDF8",x"C617",x"D679",x"E71C",x"F79D",x"FFFE",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FF3B",x"FE34",
									 x"F4A9",x"F3E3",x"F422",x"EC63",x"F483",x"FCC3",x"FCE3",x"FD04",x"FD24",x"FD44",
									 x"F564",x"FD84",x"FDA4",x"FDC6",x"FE2B",x"FEB1",x"FF35",x"FF78",x"FF59",x"FF58",
									 x"FF57",x"FF37",x"FF37",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",
									 x"FF55",x"FF55",x"FF35",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8C",x"FE8C",x"FE8B",x"FE8B",x"FE8B",
									 x"FE8A",x"FE8A",x"FE69",x"FE68",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE47",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",
									 x"FEA5",x"FEA6",x"EE05",x"BC82",x"8281",x"6120",x"58C0",x"6120",x"6960",x"6160",
									 x"6140",x"6182",x"8B6B",x"AD13",x"C618",x"CE59",x"CE38",x"CE59",x"CE79",x"CE79",
									 x"D69A",x"D69A",x"D69A",x"D69A",x"D6B9",x"D6BA",x"D6BB",x"C617",x"9CB0",x"49C4",
									 x"3120",x"4980",x"51C0",x"6221",x"7260",x"7A80",x"8AA1",x"92E2",x"A302",x"AB22",
									 x"AB42",x"B362",x"B382",x"B382",x"B383",x"B362",x"AB62",x"AB62",x"A322",x"A322",
									 x"9B02",x"9322",x"9BE2",x"B4E4",x"E6C7",x"EF67",x"FF87",x"FF66",x"FF25",x"FF05",
									 x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",
									 x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",x"FE24",x"FE04",x"FE04",x"FDC4",x"FDC4",
									 x"FDA4",x"FD64",x"FD24",x"FD03",x"FCC2",x"F483",x"EC84",x"E4CA",x"DD52",x"BDB6",
									 x"B618",x"C638",x"D6BA",x"EF5D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF9D",x"FEB8",x"F52E",x"EC26",x"F403",x"F443",
									 x"F483",x"F4A3",x"F4C3",x"FD04",x"F524",x"FD44",x"F565",x"FD85",x"FD84",x"FDA5",
									 x"FDE8",x"FE4D",x"FED2",x"FF56",x"FF79",x"FF59",x"FF78",x"FF57",x"FF36",x"FF57",
									 x"FF57",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF35",
									 x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FE8C",x"FE8C",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE69",x"FE68",
									 x"FE67",x"FE47",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE27",x"FE47",x"FE46",x"FE46",x"FE26",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE66",x"FE66",x"FE65",x"FE65",x"FE65",x"FEA5",x"FEA6",x"E5A4",x"B403",
									 x"7A01",x"5900",x"5900",x"6140",x"6960",x"6960",x"6160",x"61A2",x"8B8B",x"AD33",
									 x"C638",x"CE59",x"C638",x"CE59",x"CE79",x"CE79",x"CE79",x"CE79",x"CE79",x"D69A",
									 x"D699",x"D6DB",x"D69A",x"A533",x"83AC",x"4182",x"3940",x"49A0",x"59E0",x"6A21",
									 x"7260",x"8280",x"92C1",x"9B02",x"A302",x"AB22",x"AB42",x"B362",x"B362",x"B362",
									 x"B362",x"AB42",x"AB42",x"AB22",x"A302",x"92E2",x"9301",x"9BA1",x"B4C2",x"D625",
									 x"F767",x"FF87",x"FF66",x"FF26",x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",
									 x"FE25",x"FE24",x"FE04",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD64",x"F503",x"FCE3",
									 x"F4C2",x"F484",x"E4A7",x"D50D",x"CD94",x"BDB7",x"BE38",x"CE79",x"E71C",x"EF7D",
									 x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDF",x"FF7C",x"F633",x"ECEB",x"EC45",x"F402",x"F463",x"F483",x"F4A3",x"FCE4",
									 x"FD04",x"FD24",x"F545",x"FD65",x"FD84",x"FD85",x"FDC6",x"FE09",x"FE4D",x"FED3",
									 x"FF58",x"FF79",x"FF78",x"FF77",x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",
									 x"FF36",x"FF36",x"FF55",x"FF55",x"FF35",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8C",x"FE8C",x"FE8B",
									 x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE69",x"FE68",x"FE48",x"FE47",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE47",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",x"FE66",x"FE66",x"FE66",
									 x"FE65",x"FE85",x"FEA5",x"FE85",x"DD44",x"A363",x"6160",x"50E1",x"5920",x"6960",
									 x"6960",x"6960",x"6981",x"69E3",x"9BED",x"B554",x"C618",x"CE59",x"C638",x"C659",
									 x"CE59",x"CE79",x"CE79",x"CE79",x"CE79",x"CE79",x"D69A",x"DEDB",x"CE79",x"842F",
									 x"62A7",x"4161",x"4160",x"51C0",x"59E0",x"6A41",x"7A81",x"82A1",x"92E2",x"9B02",
									 x"A302",x"AB21",x"AB42",x"AB62",x"B342",x"B362",x"AB42",x"AB22",x"A302",x"9AE1",
									 x"92C1",x"8AE1",x"9BA1",x"C544",x"DE85",x"F786",x"FFA6",x"FF66",x"FF46",x"FF05",
									 x"FF06",x"FEE6",x"FEE6",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",
									 x"FE85",x"FE85",x"FE65",x"FE45",x"FE24",x"FE25",x"FE24",x"FE04",x"FDE4",x"FDC4",
									 x"FDA4",x"FD84",x"FD64",x"FD44",x"F4E3",x"F4C3",x"F4A3",x"ECA6",x"DCEB",x"CD51",
									 x"C5D7",x"BDF8",x"C659",x"DEDB",x"EF5D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDD",x"FEF8",x"F5D0",
									 x"F4A8",x"F402",x"F422",x"F463",x"F483",x"FCC4",x"FD04",x"F504",x"F544",x"FD65",
									 x"FD65",x"FD65",x"FD85",x"FDC6",x"FE09",x"FE8F",x"FF15",x"FF78",x"FF78",x"FF77",
									 x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF35",
									 x"FF35",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FE8C",x"FE8C",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",
									 x"FE6A",x"FE69",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE47",x"FE47",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE66",x"FE66",x"FE66",x"FE65",x"FE65",x"FE85",x"FEA6",x"FE65",
									 x"CCE4",x"92C2",x"58E0",x"50C0",x"6140",x"6960",x"6960",x"6940",x"69A2",x"7265",
									 x"A46F",x"B595",x"C617",x"C638",x"C638",x"C659",x"CE59",x"CE59",x"CE79",x"CE79",
									 x"CE79",x"CE79",x"D69A",x"DEDB",x"C637",x"6B4B",x"49E3",x"4140",x"4980",x"51C0",
									 x"6200",x"7241",x"7A81",x"82A1",x"92C2",x"9AE2",x"A301",x"AB21",x"AB22",x"AB42",
									 x"AB42",x"AB42",x"AB21",x"A301",x"9AE1",x"92C1",x"9301",x"A3E2",x"C544",x"E6A6",
									 x"F746",x"FF85",x"FF45",x"FF25",x"FF05",x"FEE5",x"FEE6",x"FEE6",x"FEE6",x"FEC5",
									 x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",
									 x"FE24",x"FE05",x"FE04",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD64",x"FD23",x"FD03",
									 x"F4C3",x"F4A3",x"EC84",x"E4E9",x"D54F",x"C5B4",x"C618",x"C638",x"D69A",x"E71C",
									 x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF7B",x"FE75",x"F50C",x"F425",x"F422",x"F442",
									 x"F483",x"F4A3",x"FCE4",x"F504",x"F524",x"FD64",x"FD64",x"FD65",x"FD85",x"FDA5",
									 x"FDC7",x"FE4B",x"FEF3",x"FF57",x"FF78",x"FF78",x"FF37",x"FF56",x"FF56",x"FF56",
									 x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF35",x"FF35",x"FF35",x"FF35",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8C",
									 x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE6A",x"FE69",x"FE68",x"FE68",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",x"FE66",
									 x"FE66",x"FE45",x"FE45",x"FE85",x"FEA6",x"F665",x"C4A3",x"8282",x"50A0",x"50C0",
									 x"6160",x"6960",x"7180",x"6140",x"69C2",x"7AC6",x"A4B0",x"BDD5",x"C617",x"C638",
									 x"C618",x"C639",x"CE59",x"CE59",x"CE79",x"CE79",x"CE79",x"CE59",x"CE79",x"D6BA",
									 x"BDD6",x"62E8",x"4181",x"4140",x"4980",x"59E0",x"6200",x"7261",x"82A1",x"8AA1",
									 x"92C1",x"A2E2",x"A301",x"AB22",x"AB22",x"A322",x"AB22",x"AB22",x"A301",x"9AE1",
									 x"92C0",x"92E1",x"A3A1",x"BD03",x"DE66",x"FF88",x"FF87",x"FF66",x"FF25",x"FF05",
									 x"FEE5",x"FEC5",x"FEC5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",
									 x"FEA5",x"FE85",x"FE85",x"FE65",x"FE45",x"FE25",x"FE04",x"FE04",x"FE04",x"FDE4",
									 x"FDC4",x"FDA4",x"FD84",x"FD43",x"FD23",x"FCE3",x"F4A3",x"F483",x"EC85",x"D50C",
									 x"D593",x"C5B6",x"BDF6",x"CE78",x"DEDB",x"EF5D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFBE",x"FEF9",x"F5B0",x"F488",x"EC03",x"F422",x"F462",x"F483",x"F4C4",x"F4E3",
									 x"F523",x"FD44",x"FD44",x"FD65",x"FD85",x"FDA5",x"FDA5",x"FDE9",x"FE90",x"FF15",
									 x"FF57",x"FF78",x"FF57",x"FF57",x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF36",
									 x"FF56",x"FF35",x"FF35",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8C",x"FE8B",x"FE8B",x"FE8B",
									 x"FE8A",x"FE8A",x"FE8A",x"FE69",x"FE68",x"FE68",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE66",x"FE45",x"FE65",x"FE85",
									 x"FE86",x"F625",x"B422",x"8222",x"50C0",x"50C0",x"6960",x"7180",x"6960",x"6140",
									 x"6A03",x"8328",x"AD32",x"BDF6",x"C617",x"C638",x"CE38",x"C639",x"CE59",x"CE59",
									 x"CE59",x"CE59",x"CE58",x"CE79",x"CE7A",x"CE79",x"A512",x"5A66",x"4140",x"4140",
									 x"51A0",x"59E0",x"6A20",x"7A61",x"82A1",x"8AA1",x"9AC2",x"A302",x"A301",x"A302",
									 x"AB22",x"A322",x"A302",x"A2E2",x"92A1",x"8AA0",x"8AE0",x"9BA1",x"BCE3",x"DE66",
									 x"F747",x"FF86",x"FF46",x"FF26",x"FF05",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",
									 x"FE45",x"FE25",x"FE04",x"FE04",x"FDE4",x"FDC4",x"FDA4",x"FDA4",x"FD63",x"FD43",
									 x"F503",x"FCE3",x"F4A3",x"EC64",x"E4C7",x"CD50",x"CDB4",x"C5F7",x"C617",x"D6BA",
									 x"E71C",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F77C",x"FE96",x"F54D",
									 x"F445",x"F423",x"F422",x"F463",x"F4C3",x"F4E3",x"FD03",x"FD24",x"FD44",x"FD64",
									 x"FD84",x"FD84",x"FDA4",x"FDA6",x"FE0B",x"FE8F",x"FF13",x"FF57",x"FF58",x"FF57",
									 x"FF57",x"FF57",x"FF56",x"FF56",x"FF56",x"FF36",x"FF36",x"FF55",x"FF35",x"FF35",
									 x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECE",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE69",
									 x"FE68",x"FE68",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE65",x"FE45",x"FE65",x"FE85",x"FE65",x"E5A5",x"A382",x"71C1",
									 x"50C0",x"58E0",x"6960",x"6981",x"6961",x"6140",x"7225",x"8B8C",x"B575",x"C617",
									 x"C618",x"BE38",x"C658",x"C658",x"CE59",x"C639",x"CE59",x"C638",x"C638",x"CE79",
									 x"D6BA",x"BDF6",x"83CD",x"51E4",x"4140",x"4980",x"59C0",x"6200",x"6A40",x"7A60",
									 x"8AA1",x"8AA1",x"92C2",x"A302",x"A2E1",x"A2E2",x"A2E2",x"A2E1",x"9AE1",x"92A1",
									 x"8A81",x"9302",x"9BE1",x"C563",x"E6A5",x"F787",x"FF86",x"FF65",x"FF25",x"FF05",
									 x"FEE5",x"FEE5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",
									 x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE04",x"FDE4",
									 x"FDE4",x"FDA4",x"FDA4",x"FD84",x"FD43",x"FD03",x"F4E4",x"F4C4",x"F484",x"E4A6",
									 x"DD2C",x"CD94",x"C5B6",x"CE18",x"CE5A",x"E71C",x"F79D",x"F7BE",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FF5A",x"FE12",x"F488",x"F403",x"F402",x"F442",
									 x"F4A3",x"F4E3",x"F4E3",x"FD04",x"FD24",x"FD44",x"FD64",x"FD84",x"F5A3",x"FDA4",
									 x"FDC7",x"FE0A",x"FEAF",x"FF54",x"FF77",x"FF58",x"FF57",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF36",x"FF36",x"FF55",x"FF35",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",
									 x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE69",x"FE68",x"FE68",x"FE67",x"FE67",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE45",x"FE65",x"FE65",
									 x"FE85",x"FE85",x"FE25",x"DD65",x"9301",x"6980",x"58E0",x"6100",x"6960",x"6960",
									 x"6960",x"6120",x"7A66",x"93CD",x"BDB6",x"C638",x"C618",x"BE18",x"C618",x"C638",
									 x"C638",x"C638",x"C638",x"C638",x"C638",x"CE7A",x"D6DA",x"B574",x"62A8",x"49A3",
									 x"4160",x"5180",x"59E1",x"6A21",x"7241",x"7A81",x"8AA1",x"8AA1",x"92C2",x"9AE1",
									 x"9AE1",x"A2E2",x"A2E2",x"9AC2",x"92A1",x"8AA1",x"9321",x"AC22",x"C564",x"E6C7",
									 x"FF68",x"FF87",x"FF46",x"FF05",x"FF05",x"FEE5",x"FEE5",x"FEE5",x"FEE5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",
									 x"FE45",x"FE45",x"FE25",x"FE05",x"FDE4",x"FDC4",x"FDC4",x"FDA4",x"F584",x"FD64",
									 x"FD23",x"F4E3",x"F4A3",x"F484",x"F486",x"DCCA",x"D56F",x"C5D5",x"BDB6",x"C618",
									 x"D69B",x"EF5D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFBD",x"FE96",x"F50C",x"E405",x"EBE2",x"F442",x"F483",x"F4C3",x"FCC3",x"FD04",
									 x"FD24",x"FD44",x"FD64",x"FD84",x"F5A4",x"FDC4",x"FDA5",x"FDC7",x"FE4B",x"FEF1",
									 x"FF56",x"FF58",x"FF57",x"FF56",x"FF56",x"FF36",x"FF36",x"FF36",x"FF36",x"FF55",
									 x"FF35",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",
									 x"FE8A",x"FE69",x"FE69",x"FE68",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE45",x"FE45",x"FE65",x"FE85",x"FE85",x"F605",x"D505",
									 x"8281",x"6120",x"58E0",x"6120",x"6960",x"6960",x"6960",x"6940",x"7AA7",x"940E",
									 x"BDB6",x"C638",x"BE18",x"BDF8",x"C618",x"C638",x"C638",x"C638",x"C618",x"C638",
									 x"CE59",x"D67A",x"D679",x"A4F2",x"5205",x"4982",x"4960",x"51A0",x"61E1",x"6A21",
									 x"7241",x"8281",x"8AA1",x"92A1",x"92A2",x"9AC1",x"9AC0",x"9AC1",x"9282",x"8A81",
									 x"8A81",x"9301",x"A421",x"C563",x"DE85",x"F767",x"FF87",x"FF46",x"FF25",x"FEE5",
									 x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",
									 x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE45",x"FE45",x"FE25",x"FE25",x"FE04",
									 x"FDC4",x"FDC4",x"FDA4",x"FD84",x"FD64",x"FD44",x"F503",x"F4E3",x"F483",x"F464",
									 x"ECA8",x"D50D",x"CD72",x"BDF7",x"BDF8",x"CE59",x"DEFC",x"EF7D",x"FFDE",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FF5B",x"FE12",x"E4AA",
									 x"EC25",x"EC23",x"F442",x"F4A3",x"FCC3",x"FCE4",x"FD04",x"FD24",x"FD44",x"FD64",
									 x"FDA4",x"FDA5",x"FD85",x"FDA6",x"FDE9",x"FE6E",x"FEF3",x"FF15",x"FF56",x"FF56",
									 x"FF56",x"FF36",x"FF36",x"FF56",x"FF36",x"FF35",x"FF35",x"FF35",x"FF35",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF33",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FF12",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",
									 x"FECD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE69",x"FE68",
									 x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE45",x"FE65",x"FE85",x"FE85",x"EDC4",x"C464",x"71E0",x"58E0",x"6100",x"6940",
									 x"7160",x"7180",x"7160",x"7181",x"82C7",x"9C4F",x"B5B6",x"C618",x"BE18",x"BDF8",
									 x"C5F8",x"C618",x"C638",x"C638",x"BE18",x"C618",x"CE59",x"CE18",x"B594",x"8BED",
									 x"4182",x"4960",x"4980",x"59C1",x"6A01",x"7221",x"7A41",x"8261",x"8A81",x"9281",
									 x"92A1",x"9AA1",x"92A0",x"9281",x"8A60",x"8AA0",x"9341",x"B4A4",x"DE46",x"F726",
									 x"FF66",x"FF66",x"FF26",x"FF05",x"FF05",x"FEE5",x"FEE5",x"FEC6",x"FEC5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",
									 x"FE65",x"FE45",x"FE25",x"FE25",x"FE05",x"FDE5",x"FDC4",x"FDC4",x"FDA4",x"FD64",
									 x"FD44",x"FD24",x"FCE3",x"F4C2",x"F482",x"EC65",x"DD0C",x"CD71",x"C5D4",x"BE18",
									 x"C659",x"D6BB",x"E73D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"FEB7",x"ED4F",x"F4A8",x"EC43",x"EC22",x"F462",
									 x"F4A3",x"F4C3",x"FCE4",x"FD04",x"FD24",x"FD44",x"FD85",x"FDA5",x"FD65",x"FD85",
									 x"FDA6",x"F60A",x"FE8F",x"FED2",x"FF35",x"FF57",x"FF57",x"FF56",x"FF56",x"FF36",
									 x"FF36",x"FF35",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF33",
									 x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FEAD",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8A",
									 x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE69",x"FE68",x"FE68",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE45",x"FE45",x"FE65",x"FE85",x"FE65",
									 x"E584",x"ABC2",x"6140",x"50A0",x"6101",x"6960",x"7180",x"7180",x"7180",x"79E2",
									 x"8B29",x"A4B1",x"B5B6",x"BE18",x"BDF8",x"BDD8",x"C5F8",x"C5F7",x"C617",x"C618",
									 x"C659",x"C659",x"CE39",x"AD13",x"7BAC",x"5A66",x"4161",x"51A0",x"51C0",x"59E0",
									 x"7201",x"7A21",x"8241",x"8A61",x"8A61",x"9282",x"8A61",x"8A60",x"8A40",x"8A61",
									 x"9302",x"A3C1",x"BCE3",x"E687",x"F747",x"FF86",x"FF45",x"FF06",x"FEE6",x"FEE5",
									 x"FEE5",x"FEC5",x"FEC5",x"FEC6",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",
									 x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE05",
									 x"FDE5",x"FDE5",x"FDC4",x"FDA4",x"FD84",x"FD64",x"FD24",x"FD04",x"F4C3",x"F482",
									 x"F484",x"E4A9",x"D550",x"CDD5",x"C5F6",x"C659",x"D6BA",x"E71B",x"F79E",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",
									 x"FF3B",x"F613",x"F52C",x"EC24",x"EC22",x"F442",x"F483",x"F4C3",x"FCE4",x"FD04",
									 x"FD24",x"FD44",x"FD64",x"FD84",x"FD65",x"FD85",x"FDA5",x"FDE6",x"FE2A",x"FE8F",
									 x"FF14",x"FF58",x"FF58",x"FF56",x"FF55",x"FF36",x"FF36",x"FF35",x"FF35",x"FF35",
									 x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF33",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",
									 x"FE69",x"FE68",x"FE68",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE26",x"FE45",x"FE65",x"FE85",x"FE45",x"D524",x"A362",x"6120",x"5080",
									 x"6121",x"7180",x"7180",x"7180",x"7980",x"7A02",x"936A",x"A4B1",x"B5D7",x"BE18",
									 x"B5F8",x"BDF8",x"BE18",x"C618",x"C638",x"C639",x"C659",x"C639",x"BDD6",x"942F",
									 x"6287",x"51E3",x"4160",x"51A0",x"59C0",x"6201",x"7221",x"7A21",x"8261",x"8A81",
									 x"8A62",x"8A42",x"8A41",x"8240",x"8241",x"8AC2",x"9BC2",x"B4C2",x"D624",x"FF88",
									 x"FFA7",x"FF66",x"FF25",x"FEE5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",
									 x"FE65",x"FE45",x"FE45",x"FE25",x"FE05",x"FE04",x"FDE5",x"FDC4",x"FDA4",x"FD84",
									 x"FD84",x"F544",x"FD03",x"FCC3",x"F483",x"F483",x"EC87",x"DCED",x"CD95",x"BDF7",
									 x"BE17",x"CE79",x"DEDB",x"EF5C",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"F6F8",x"FE12",x"EC88",
									 x"EC24",x"F402",x"F442",x"F483",x"F4C3",x"F4E4",x"F504",x"FD24",x"FD44",x"FD64",
									 x"FD64",x"FD85",x"F584",x"FDA5",x"FDE6",x"FE2A",x"FEB0",x"FF35",x"FF57",x"FF56",
									 x"FF55",x"FF35",x"FF35",x"FF35",x"FF35",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FEF2",x"FEF2",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",
									 x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE69",x"FE68",x"FE67",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE26",x"FE25",x"FE65",
									 x"FE85",x"F605",x"C4A3",x"92E3",x"5900",x"50A0",x"6940",x"7161",x"7180",x"7980",
									 x"7980",x"7A03",x"936A",x"A4B1",x"B5D7",x"BE39",x"B618",x"BE38",x"BE39",x"BE39",
									 x"BE18",x"BDF7",x"B5B6",x"AD34",x"942E",x"6267",x"4982",x"4981",x"5180",x"59C0",
									 x"61C0",x"6A01",x"7221",x"7A41",x"8241",x"8261",x"8221",x"8201",x"8200",x"8A61",
									 x"8B02",x"A423",x"D5E6",x"EF06",x"F786",x"FFA6",x"F725",x"FF05",x"FEE5",x"FEC5",
									 x"FEA5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",
									 x"FE05",x"FDE5",x"FDC4",x"FDA4",x"FD84",x"FD64",x"F564",x"F523",x"FCE3",x"FCA3",
									 x"F484",x"ECA5",x"DCCA",x"D551",x"C5B6",x"BDF7",x"BE58",x"D6BA",x"E71C",x"EF7D",
									 x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FF9D",x"FF18",x"ED8F",x"E467",x"EC03",x"EC22",x"F462",
									 x"F483",x"F4C3",x"F4E3",x"F504",x"F524",x"FD44",x"FD64",x"FD64",x"FD84",x"F584",
									 x"F5A5",x"F5E7",x"FE4B",x"FEB0",x"FF14",x"FF55",x"FF76",x"FF55",x"FF35",x"FF35",
									 x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF12",x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",
									 x"FE8A",x"FE8A",x"FE69",x"FE68",x"FE68",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE45",x"FE85",x"FE66",x"E5A4",x"ABE2",x"7A21",
									 x"58E0",x"58E0",x"6940",x"7181",x"7981",x"7980",x"7980",x"79C2",x"8AE8",x"9C0E",
									 x"B554",x"BDD6",x"B5B6",x"B5D6",x"B5B6",x"B575",x"AD12",x"9C90",x"83AC",x"7B4A",
									 x"5A04",x"4140",x"4140",x"4960",x"59C0",x"6200",x"61E0",x"6A01",x"7A20",x"7A20",
									 x"7A00",x"7A21",x"8221",x"8241",x"8AE0",x"AC22",x"C524",x"DE46",x"F747",x"FFA7",
									 x"FF66",x"FF05",x"FF05",x"FEE5",x"FEE6",x"FEC6",x"FEA5",x"FEA5",x"FEA5",x"FEA5",
									 x"FEA5",x"FEA5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",
									 x"FE65",x"FE65",x"FE45",x"FE25",x"FE25",x"FE05",x"FE05",x"FDE4",x"FDC4",x"FDA4",
									 x"FD64",x"FD44",x"F544",x"F502",x"FCC2",x"F483",x"EC85",x"E4C9",x"D52D",x"CDB3",
									 x"BDD6",x"BE18",x"CE99",x"E73C",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",
									 x"FF9D",x"F676",x"E50C",x"EC45",x"F422",x"F442",x"F462",x"F4A3",x"F4E3",x"F504",
									 x"F504",x"FD44",x"FD65",x"FD65",x"FD84",x"FD85",x"F5A5",x"F5C5",x"FDE8",x"FE2B",
									 x"FE90",x"FF14",x"FF56",x"FF56",x"FF36",x"FF35",x"FF35",x"FF34",x"FF34",x"FF34",
									 x"FF34",x"FF34",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",
									 x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FE8C",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",
									 x"FE68",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE65",x"FE85",x"FE46",x"D524",x"9B41",x"6180",x"50C0",x"5900",x"6940",x"7181",
									 x"7981",x"7980",x"7980",x"7180",x"8265",x"9349",x"A46F",x"ACF1",x"ACF1",x"A4D1",
									 x"9C90",x"942F",x"93AB",x"7AE8",x"51E4",x"4981",x"4140",x"4960",x"5180",x"51A0",
									 x"61C0",x"61E0",x"69E0",x"7201",x"7A00",x"79E0",x"71E0",x"7A00",x"82A1",x"9341",
									 x"AC81",x"DE25",x"EEC6",x"F766",x"FF66",x"FF45",x"FF05",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA6",x"FEA6",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",
									 x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",x"FE45",x"FE25",
									 x"FE25",x"FE05",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD64",x"FD43",x"F503",x"F4C2",
									 x"FCA2",x"EC84",x"E4C8",x"DD2E",x"CD91",x"C5F5",x"BE18",x"CE59",x"DEBA",x"EF7D",
									 x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FF1A",x"EDB0",x"F4A9",
									 x"EC24",x"EC23",x"F442",x"F483",x"F4C3",x"F4E4",x"F504",x"FD24",x"FD45",x"FD65",
									 x"FD65",x"FD85",x"FDA6",x"F5A6",x"FDA6",x"FDE8",x"FE2C",x"FEB1",x"FF15",x"FF36",
									 x"FF36",x"FF36",x"FF16",x"FF15",x"FF15",x"FF35",x"FF34",x"FF34",x"FF34",x"FF34",
									 x"FF14",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FEF2",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",
									 x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE69",x"FE68",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE27",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE47",x"FE46",
									 x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE65",x"FE85",x"F627",x"CCC5",
									 x"8281",x"50E0",x"50A0",x"6120",x"7160",x"7160",x"7981",x"79A1",x"79A0",x"79A1",
									 x"81E2",x"8A64",x"8B08",x"9389",x"938A",x"8B6A",x"7AE8",x"7286",x"6A25",x"59E3",
									 x"4981",x"4960",x"4960",x"51A1",x"59A1",x"61A1",x"61C1",x"61A0",x"69C0",x"61A0",
									 x"71C1",x"71E1",x"7A20",x"8AE1",x"A422",x"BCE3",x"D624",x"EF06",x"F746",x"FF66",
									 x"FF46",x"FEE5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA6",x"FEA6",x"FEC5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",
									 x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE25",x"FE05",x"FE05",x"FDE4",x"FDC4",
									 x"FD84",x"FD64",x"FD44",x"FD23",x"F4E3",x"F4A2",x"F483",x"E486",x"DCEB",x"D592",
									 x"C5B4",x"BDF6",x"C659",x"D69A",x"E6FB",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FF9D",x"FE96",x"F5AF",x"F4A8",x"EC04",x"F423",x"F463",
									 x"F483",x"F4C3",x"F4E4",x"FD04",x"FD24",x"FD45",x"FD65",x"FD85",x"FDA6",x"FDA6",
									 x"FDA5",x"FDA6",x"FDC8",x"FE2C",x"FEB0",x"FF14",x"FF35",x"FF36",x"FF36",x"FF15",
									 x"FF15",x"FF35",x"FF15",x"FF34",x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",
									 x"FF13",x"FF12",x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE89",
									 x"FE89",x"FE89",x"FE69",x"FE68",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE47",
									 x"FE47",x"FE47",x"FE46",x"FE46",x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",
									 x"FE45",x"FE45",x"FE65",x"FE86",x"EDC6",x"B403",x"7201",x"4060",x"50C1",x"6140",
									 x"7160",x"7160",x"79A1",x"79A1",x"79A1",x"79A0",x"7980",x"79A0",x"79C1",x"7A01",
									 x"71E2",x"61A1",x"5960",x"5100",x"4920",x"5140",x"51A1",x"59C1",x"59A1",x"61C2",
									 x"61A1",x"61A1",x"69A1",x"69A0",x"69C0",x"69C0",x"7201",x"82A1",x"9BA1",x"BCE3",
									 x"DE25",x"EEE6",x"FF87",x"FF87",x"FF46",x"FF05",x"FEC5",x"FEA5",x"FEA5",x"FEA5",
									 x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",
									 x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE25",
									 x"FE25",x"FE05",x"FE05",x"FDE4",x"FDC4",x"FDA3",x"FD84",x"FD44",x"F504",x"F4E4",
									 x"F4A3",x"F463",x"EC65",x"DCCA",x"D52F",x"CDD5",x"C5D6",x"C617",x"D69A",x"DEFB",
									 x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",
									 x"FF5B",x"FE96",x"FD4D",x"EC46",x"EC03",x"F422",x"F442",x"F4A3",x"F4C3",x"F4E4",
									 x"FD04",x"FD24",x"FD44",x"FD65",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDE7",
									 x"FE4B",x"FEB0",x"FF13",x"FF55",x"FF56",x"FF34",x"FF34",x"FF15",x"FF15",x"FF14",
									 x"FF34",x"FF34",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",x"FEF2",x"FEF2",
									 x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8B",
									 x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE8A",x"FE8A",x"FE69",x"FE68",
									 x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",
									 x"FE47",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE46",x"FE45",x"FE65",x"FE66",
									 x"DD65",x"9B62",x"6180",x"3840",x"50C0",x"6140",x"6960",x"7160",x"79A0",x"79A0",
									 x"79C0",x"81E0",x"79C0",x"81C0",x"79C0",x"79C0",x"71A0",x"69A0",x"69A0",x"6160",
									 x"6160",x"5980",x"61A0",x"61A0",x"61A0",x"61A0",x"6181",x"6160",x"6180",x"71E0",
									 x"7220",x"8AC1",x"9BC2",x"B4C3",x"D5E4",x"EEC5",x"F745",x"FF45",x"FF25",x"FF05",
									 x"FEE5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEC5",x"FEC5",
									 x"FEC5",x"FEC5",x"FEC5",x"FEC5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",
									 x"FE65",x"FE65",x"FE65",x"FE45",x"FE25",x"FE25",x"FE05",x"FE05",x"FDE4",x"FDC4",
									 x"FDA4",x"FD83",x"FD63",x"F524",x"F4E4",x"F4C3",x"F482",x"F484",x"EC87",x"DD0D",
									 x"CD92",x"C5F6",x"C5F7",x"CE59",x"E6FC",x"EF5D",x"F7BE",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FF9D",x"FF3A",x"F613",x"E4CA",
									 x"E404",x"F402",x"FC22",x"FCA2",x"F4C3",x"F4C4",x"FD04",x"FD24",x"FD44",x"FD64",
									 x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FE07",x"FE6C",x"FED1",x"FF15",
									 x"FF36",x"FF15",x"FF14",x"FF15",x"FF14",x"FF34",x"FF14",x"FF14",x"FF14",x"FF13",
									 x"FF13",x"FF13",x"FF12",x"FF12",x"FF11",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",
									 x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE69",x"FE69",x"FE68",x"FE67",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE27",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE47",x"FE46",x"FE26",x"FE26",
									 x"FE26",x"FE46",x"FE46",x"FE46",x"FE65",x"FE65",x"D504",x"92E2",x"5961",x"4080",
									 x"50E0",x"6140",x"6940",x"7140",x"7981",x"7980",x"79A0",x"81C0",x"79C0",x"79A0",
									 x"71A0",x"71A0",x"71A0",x"69C0",x"69C0",x"69C0",x"69C0",x"61A0",x"6181",x"6181",
									 x"6180",x"6180",x"6981",x"6981",x"71E0",x"82C1",x"9361",x"AC62",x"C582",x"D643",
									 x"EEE5",x"FF66",x"FF66",x"FF45",x"FEE5",x"FEC5",x"FEC5",x"FEA5",x"FE84",x"FE85",
									 x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",
									 x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",
									 x"FE25",x"FE05",x"FDE5",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD64",x"FD43",x"F523",
									 x"F4E3",x"F4A2",x"EC82",x"ECC6",x"DCEB",x"CD71",x"C5F5",x"BDF7",x"C618",x"D6BA",
									 x"E73C",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFDE",x"FFBC",x"FF19",x"EDD1",x"E489",x"F424",x"F403",x"F463",
									 x"F483",x"F4A3",x"F4E4",x"F504",x"F524",x"FD44",x"FD64",x"F564",x"FDA5",x"FDC5",
									 x"FDA5",x"FDA5",x"FDC6",x"FDE9",x"FE4C",x"FEB0",x"FEF3",x"FF35",x"FF35",x"FF34",
									 x"FF34",x"FF34",x"FF33",x"FF33",x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FF12",
									 x"FF12",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",
									 x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE8A",
									 x"FE69",x"FE69",x"FE68",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE47",x"FE47",x"FE47",
									 x"FE46",x"FE46",x"FE47",x"FE46",x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE46",
									 x"FE65",x"F645",x"C4A4",x"8281",x"5121",x"4060",x"50C1",x"5921",x"6940",x"6941",
									 x"7961",x"7981",x"7981",x"79A1",x"79A1",x"79A1",x"79C1",x"79C0",x"79C0",x"71C1",
									 x"71C1",x"69C1",x"69A0",x"6160",x"5940",x"5100",x"5940",x"61A0",x"7260",x"82E0",
									 x"9BC2",x"BCE4",x"CDC4",x"EEA6",x"FF27",x"FF47",x"FF26",x"FF05",x"FEE5",x"FEC4",
									 x"FEA5",x"FE85",x"FE84",x"FEA5",x"FE85",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",
									 x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE25",x"FE04",x"FDE4",x"FDE4",x"FDC4",
									 x"FDC4",x"FDA4",x"FD64",x"F543",x"FD22",x"FCE3",x"F483",x"F463",x"E4A6",x"DCEA",
									 x"DD50",x"CDB5",x"C5F7",x"C638",x"D69A",x"E71C",x"F79E",x"F7BE",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",
									 x"FFBE",x"F6D9",x"F58F",x"FCA9",x"EBE4",x"F403",x"F442",x"F483",x"F4A3",x"F4C4",
									 x"F4E3",x"FD24",x"FD44",x"F544",x"FD65",x"FD85",x"FDA5",x"FDA5",x"FD85",x"FD85",
									 x"FDE7",x"F64A",x"FE8E",x"FED2",x"FEF4",x"FF15",x"FF35",x"FF34",x"FF34",x"FF13",
									 x"FF13",x"FF13",x"FF13",x"FF13",x"FF12",x"FEF2",x"FF12",x"FEF2",x"FEF1",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8B",x"FE8B",x"FE8B",
									 x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE8A",x"FE8A",x"FE69",x"FE69",x"FE68",x"FE67",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE27",x"FE47",x"FE47",x"FE47",x"FE46",x"FE46",x"FE47",x"FE46",
									 x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE46",x"FE66",x"F646",x"C4A4",x"7A60",
									 x"5100",x"4060",x"50E1",x"5920",x"6140",x"6940",x"7160",x"7980",x"7980",x"79A0",
									 x"79A0",x"79A0",x"7961",x"7140",x"6940",x"6120",x"6120",x"6120",x"6160",x"69C1",
									 x"7222",x"7A61",x"8B02",x"A3E4",x"B4C3",x"C564",x"E666",x"EEE6",x"F726",x"F745",
									 x"FF26",x"FF06",x"FEE5",x"FEA5",x"FE85",x"FE85",x"FEA5",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FEA5",x"FE85",x"FE85",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",x"FEA5",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",x"FE45",x"FE25",x"FE25",
									 x"FE25",x"FE04",x"FDE4",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD64",x"F544",x"F523",
									 x"F4E2",x"FC83",x"FC44",x"F465",x"DCCA",x"D570",x"CDB5",x"C5D7",x"CE39",x"D6BA",
									 x"DEFB",x"EF7D",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F75B",x"FE54",x"FD2D",
									 x"F427",x"F403",x"F423",x"F463",x"F4A3",x"F4C4",x"F4E3",x"FD04",x"FD24",x"FD44",
									 x"FD65",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FD84",x"FDC4",x"FE06",x"FE4A",x"FE8F",
									 x"FED2",x"FF14",x"FF15",x"FF35",x"FF35",x"FF14",x"FF14",x"FF13",x"FF13",x"FF13",
									 x"FEF2",x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FE8C",x"FEAB",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE89",
									 x"FE89",x"FE8A",x"FE69",x"FE69",x"FE68",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE45",x"FE46",x"FE45",x"FE46",x"CCE4",x"82A0",x"5101",x"3840",x"48A1",x"50E1",
									 x"5900",x"6121",x"6921",x"6921",x"7141",x"7161",x"7160",x"7160",x"7141",x"7141",
									 x"6941",x"6961",x"6960",x"6980",x"71E0",x"8282",x"9363",x"A3E2",x"B4A2",x"CDA4",
									 x"E645",x"EEC6",x"FF47",x"FF67",x"FF46",x"F704",x"F6A4",x"FEA5",x"FE85",x"FE85",
									 x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FEA5",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE45",x"FE25",x"FE25",x"FE25",x"FE05",x"FE05",x"FDE4",x"FDC4",
									 x"FDA4",x"FD84",x"FD84",x"FD44",x"F523",x"F503",x"FCC2",x"F463",x"F445",x"E4A8",
									 x"D52D",x"CDB3",x"C5F7",x"C5F7",x"CE79",x"DEFB",x"E73C",x"F7BE",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"FF39",x"FE34",x"ECEC",x"EC25",x"EC02",x"EC22",
									 x"F463",x"FCA4",x"FCC3",x"FCE4",x"FD04",x"FD24",x"FD45",x"FD65",x"FD65",x"FD85",
									 x"FDA5",x"FDA5",x"FDA4",x"FDC5",x"FE07",x"FE2B",x"FE6D",x"FED0",x"FEF2",x"FF34",
									 x"FF35",x"FF14",x"FF14",x"FF13",x"FF13",x"FF13",x"FEF2",x"FEF2",x"FEF2",x"FEF1",
									 x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAB",
									 x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE89",x"FE69",x"FE69",
									 x"FE68",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE26",x"FE45",x"FE65",
									 x"DD65",x"9B42",x"6161",x"3820",x"3820",x"4061",x"4880",x"50A1",x"58A0",x"58A0",
									 x"58A0",x"58E0",x"6100",x"6120",x"7180",x"79E1",x"7A20",x"8260",x"8AE1",x"9342",
									 x"A3C1",x"B463",x"CD65",x"DDE5",x"E665",x"EEA5",x"F6E6",x"FEE6",x"FEE5",x"FEE5",
									 x"FEC5",x"FEA5",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE64",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE25",
									 x"FE25",x"FE05",x"FE05",x"FDE4",x"FDC4",x"FDA4",x"FDA4",x"FD64",x"F563",x"F523",
									 x"FD03",x"FCC2",x"F482",x"EC65",x"E488",x"DD0D",x"CDB1",x"C5F5",x"BDF7",x"C638",
									 x"D6BA",x"E73C",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",
									 x"FFDE",x"FF3B",x"FE14",x"F4EB",x"F465",x"F422",x"F442",x"F463",x"F483",x"F4C3",
									 x"FCE4",x"FD04",x"FD24",x"FD44",x"FD64",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",
									 x"FDC6",x"FDC7",x"FDE8",x"FE4B",x"FEAE",x"FEF1",x"FF13",x"FF14",x"FF14",x"FF14",
									 x"FF13",x"FEF3",x"FEF2",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FEF1",
									 x"FEF1",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAB",x"FE8B",x"FE8B",x"FE8A",x"FE8A",
									 x"FE8A",x"FE89",x"FE89",x"FE89",x"FE69",x"FE69",x"FE68",x"FE68",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE46",x"FE46",x"FE45",x"FE65",x"EDE6",x"C484",x"8AE2",x"61A0",
									 x"5100",x"5120",x"5940",x"6140",x"6160",x"6981",x"69A1",x"7201",x"7A21",x"8A81",
									 x"9B22",x"A3A3",x"AC22",x"BCC3",x"CD64",x"D5E4",x"E624",x"EE85",x"F6C6",x"FF06",
									 x"FF26",x"FF06",x"FEC5",x"FEC4",x"FE84",x"FE64",x"FE45",x"FE46",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE85",x"FE84",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",
									 x"FE65",x"FE45",x"FE45",x"FE25",x"FE25",x"FE25",x"FE05",x"FDE5",x"FDE4",x"FDC4",
									 x"FDA4",x"FD84",x"FD84",x"F543",x"F543",x"F503",x"FCC2",x"FC82",x"F483",x"E4A7",
									 x"DCEC",x"D572",x"CDF5",x"C617",x"CE59",x"D69A",x"E73C",x"F7BE",x"FFDF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FEF9",x"F5D1",
									 x"ECCA",x"EC04",x"F3E2",x"FC42",x"F463",x"F4A4",x"F4C4",x"F4E4",x"F524",x"FD24",
									 x"FD44",x"FD64",x"FD65",x"FD84",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC6",x"FDE7",
									 x"FE49",x"FE8C",x"FED0",x"FF13",x"FF14",x"FF14",x"FF13",x"FF13",x"FEF2",x"FEF2",
									 x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FED1",x"FEF0",x"FED0",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FE8C",x"FEAB",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE89",
									 x"FE89",x"FE69",x"FE68",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE45",
									 x"FE45",x"FE45",x"FE46",x"EDE6",x"CCE5",x"AC03",x"9322",x"82C1",x"8AE2",x"8B02",
									 x"9B42",x"A383",x"ABE3",x"B443",x"BC83",x"CCE4",x"D564",x"DDC5",x"E625",x"F6A5",
									 x"F6E5",x"FF25",x"FF25",x"FF05",x"FEE5",x"FEA5",x"FEA5",x"FE85",x"FE64",x"FE64",
									 x"FE44",x"FE65",x"FE45",x"FE45",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE85",x"FE85",x"FE65",x"FE65",x"FE45",x"FE45",x"FE25",x"FE25",
									 x"FE04",x"FE04",x"FDE4",x"FDC4",x"FDC4",x"FDA4",x"FD84",x"FD84",x"FD44",x"FD04",
									 x"FD03",x"F4E3",x"F482",x"F462",x"E485",x"DCEB",x"D551",x"C5B5",x"C5F7",x"C638",
									 x"D6BA",x"DEFC",x"F77E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FF7C",x"FE97",x"F5B1",x"E489",x"EC04",x"F423",
									 x"F443",x"F4A4",x"F4A3",x"F4C3",x"F4E4",x"F504",x"FD24",x"FD44",x"FD64",x"FD64",
									 x"FD85",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDC6",x"FDE7",x"FE29",x"FE6C",x"FECF",
									 x"FF11",x"FEF3",x"FF13",x"FF13",x"FEF3",x"FEF3",x"FEF2",x"FEF2",x"FEF1",x"FEF1",
									 x"FEF1",x"FEF1",x"FED1",x"FEF0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FEAB",x"FE8B",x"FE8B",
									 x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE89",x"FE89",x"FE69",x"FE68",x"FE68",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",x"FE46",x"FE45",x"FE45",x"FE46",x"FE26",
									 x"E5C5",x"D544",x"C4A3",x"BC63",x"BC63",x"BC83",x"C4C3",x"CD24",x"D544",x"DDA4",
									 x"E5C4",x"E5E4",x"EE44",x"F665",x"F685",x"FEC5",x"FEE5",x"FEE5",x"FEE5",x"FEC5",
									 x"FEA5",x"FE85",x"FE65",x"FE45",x"FE65",x"FE44",x"FE44",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",x"FE05",x"FE04",x"FDE4",x"FDC4",x"FDC4",
									 x"FDA4",x"FD84",x"F584",x"F564",x"FD23",x"FCE3",x"FCC3",x"F4A3",x"F463",x"EC85",
									 x"DCC9",x"D52F",x"D594",x"C5D6",x"C617",x"CE9A",x"DF1C",x"EF5D",x"FFBE",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDE",x"FF5C",x"F6B8",x"ED90",x"EC68",x"F404",x"F402",x"F463",x"F483",x"F4A3",
									 x"F4C4",x"FD04",x"F504",x"FD24",x"FD44",x"FD64",x"FD64",x"FD85",x"FDA5",x"FDA5",
									 x"FDC5",x"FDA5",x"FDC5",x"FDE6",x"FE28",x"FE6B",x"FEAC",x"FECF",x"FEF1",x"FEF3",
									 x"FF14",x"FF13",x"FEF2",x"FEF2",x"FEF1",x"FEF1",x"FEF1",x"FEF1",x"FED1",x"FEF0",
									 x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",
									 x"FECE",x"FECD",x"FECD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FE8C",x"FEAB",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE89",
									 x"FE89",x"FE89",x"FE89",x"FE69",x"FE68",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE25",x"FE45",x"FE46",x"FE46",x"FE65",x"FE65",x"FE46",x"F626",
									 x"F625",x"F645",x"F686",x"FEA6",x"FEC6",x"FEC6",x"FEC6",x"FEC5",x"FEC5",x"FEA4",
									 x"FE84",x"FE84",x"FE84",x"FE64",x"FE44",x"FE44",x"FE45",x"FE44",x"FE45",x"FE45",
									 x"FE45",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",x"FE85",x"FE85",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",
									 x"FE05",x"FE05",x"FDE4",x"FDE4",x"FDC4",x"FDA4",x"FD84",x"FD84",x"F543",x"F523",
									 x"FD03",x"FCC3",x"F482",x"F463",x"EC86",x"E4EA",x"D52E",x"CDB3",x"C5D6",x"CE17",
									 x"CE79",x"DF1B",x"EF7E",x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FF9D",x"FEB7",
									 x"FD6E",x"F467",x"F404",x"F402",x"F442",x"F462",x"F4A3",x"F4C4",x"F4E4",x"F504",
									 x"FD24",x"FD44",x"FD44",x"FD65",x"FD85",x"FDA5",x"FDA5",x"FDC5",x"FDA5",x"FDC5",
									 x"FDE6",x"FE07",x"FE49",x"FE8B",x"FEAE",x"FED1",x"FEF3",x"FF13",x"FEF2",x"FEF2",
									 x"FEF2",x"FEF1",x"FED1",x"FED1",x"FED1",x"FEF0",x"FEF0",x"FED0",x"FED0",x"FECF",
									 x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FEAD",x"FEAD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8B",
									 x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE89",x"FE89",x"FE69",
									 x"FE68",x"FE68",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE45",x"FE25",
									 x"FE25",x"FE25",x"FE44",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE85",
									 x"FE85",x"FE85",x"FE85",x"FE85",x"FE85",x"FE64",x"FE65",x"FE45",x"FE45",x"FE25",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE64",x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",x"FE05",x"FE05",x"FDE4",x"FDC4",x"FDC4",
									 x"FDA4",x"FD84",x"FD84",x"FD64",x"F523",x"F502",x"FCE3",x"F4A3",x"F483",x"EC85",
									 x"E4CA",x"DD4F",x"CDB3",x"C5D6",x"C618",x"CE79",x"DEFB",x"EF7D",x"F7DF",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FF5B",x"F613",x"ED0C",x"EC67",x"EC03",
									 x"F422",x"F442",x"F483",x"F4A3",x"F4E3",x"FD04",x"FD24",x"FD24",x"FD44",x"FD65",
									 x"FD65",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FE06",x"FE07",x"FE28",
									 x"FE6A",x"FE8D",x"FEAF",x"FED1",x"FEF1",x"FEF1",x"FEF2",x"FEF2",x"FEF2",x"FED1",
									 x"FED0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",
									 x"FECE",x"FECE",x"FECE",x"FEAD",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",
									 x"FE8A",x"FE89",x"FE89",x"FE89",x"FE69",x"FE69",x"FE68",x"FE48",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE46",x"FE25",x"FE25",x"FE25",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE65",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",x"FE05",
									 x"FE05",x"FE05",x"FDE5",x"FDC4",x"FDC4",x"FDA4",x"FD84",x"FD63",x"FD44",x"FD23",
									 x"FD03",x"FCC2",x"F4A3",x"F484",x"EC65",x"E4A8",x"D50E",x"CD93",x"C5F5",x"C617",
									 x"CE59",x"D6BA",x"E73C",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFDE",x"FF19",x"F634",x"ED4E",x"EC66",x"EC23",x"F422",x"F463",x"F483",
									 x"F4A3",x"F4E3",x"FD04",x"FD04",x"FD24",x"FD44",x"FD45",x"FD65",x"FD85",x"FDA6",
									 x"FDA6",x"FDC5",x"FDC6",x"FDC6",x"FDC6",x"FDE6",x"FE07",x"FE49",x"FE6B",x"FE8E",
									 x"FEB0",x"FED1",x"FED1",x"FEF2",x"FED1",x"FED1",x"FED0",x"FED0",x"FED0",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECE",x"FEAD",
									 x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE89",
									 x"FE89",x"FE69",x"FE68",x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE45",x"FE45",
									 x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",x"FE25",x"FE45",x"FE45",x"FE44",
									 x"FE64",x"FE64",x"FE65",x"FE65",x"FE65",x"FE64",x"FE64",x"FE64",x"FE44",x"FE64",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE25",x"FE24",x"FE04",x"FE04",x"FDE4",x"FDE4",x"FDE4",x"FDC4",
									 x"FDA4",x"FD84",x"FD64",x"FD43",x"FD23",x"FCE3",x"FCC2",x"F4A2",x"F483",x"EC85",
									 x"E4A7",x"DD0C",x"D572",x"C5D6",x"BE17",x"CE58",x"DEDA",x"E73C",x"F79E",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FFBC",x"FF7B",
									 x"FE96",x"F54D",x"EC87",x"EC25",x"F423",x"F443",x"F483",x"F4A3",x"F4C3",x"FCE3",
									 x"FD04",x"FD24",x"FD44",x"FD64",x"FD65",x"FD85",x"FDA5",x"FDA5",x"FDC5",x"FDC5",
									 x"FDC5",x"FDC5",x"FDC5",x"FDE6",x"FE08",x"FE29",x"FE6B",x"FE8D",x"FEAE",x"FEB0",
									 x"FED1",x"FED1",x"FEF0",x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECF",
									 x"FECF",x"FECE",x"FECE",x"FEAE",x"FEAE",x"FECD",x"FEAD",x"FEAD",x"FEAD",x"FEAC",
									 x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",
									 x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE89",x"FE89",x"FE68",x"FE68",x"FE67",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE65",x"FE65",
									 x"FE65",x"FE45",x"FE45",x"FE45",x"FE64",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE85",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",x"FE24",x"FE04",
									 x"FE04",x"FDE4",x"FDE4",x"FDC4",x"FDA4",x"FDA3",x"FD83",x"FD64",x"FD44",x"FD24",
									 x"FD03",x"FCC3",x"F483",x"F483",x"ECA5",x"E4C9",x"D52D",x"D592",x"CDD5",x"C617",
									 x"C659",x"DEDB",x"EF5D",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",x"FFDE",x"FF5C",x"FE75",x"ED4D",x"ECA9",
									 x"F424",x"F402",x"EC22",x"F462",x"FCA3",x"F4C3",x"FD04",x"F504",x"F524",x"FD64",
									 x"FD64",x"FD64",x"FD85",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDA5",x"FDC5",x"FDC5",
									 x"FDE6",x"FDE7",x"FE08",x"FE2A",x"FE4B",x"FE6C",x"FEAE",x"FECF",x"FED0",x"FED0",
									 x"FED0",x"FED0",x"FED0",x"FED0",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FECD",
									 x"FEAD",x"FEAD",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",
									 x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",
									 x"FE8A",x"FE89",x"FE69",x"FE68",x"FE68",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE44",x"FE44",
									 x"FE24",x"FE25",x"FE25",x"FE05",x"FE04",x"FE04",x"FDE4",x"FDE4",x"FDC4",x"FDA4",
									 x"FD84",x"FD83",x"FD63",x"FD23",x"F503",x"FCE3",x"FCC2",x"FC82",x"F463",x"EC85",
									 x"E4E9",x"DD4E",x"D592",x"CDF5",x"CE37",x"CE79",x"D6DB",x"E75D",x"F7BE",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFDF",x"FF5B",x"F675",x"F5B0",x"EC88",x"F403",x"F402",x"F422",
									 x"F463",x"F4C3",x"F4E4",x"F4E4",x"F504",x"F524",x"FD44",x"FD44",x"FD64",x"FD65",
									 x"FD85",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDC5",x"FDE6",x"FDE6",x"FDE6",x"FE07",
									 x"FE27",x"FE48",x"FE6A",x"FE8C",x"FE8E",x"FEAF",x"FEAF",x"FED0",x"FEF1",x"FED0",
									 x"FED0",x"FECF",x"FECF",x"FECE",x"FECE",x"FECE",x"FEAE",x"FEAE",x"FEAD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8C",x"FE8B",
									 x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE6A",x"FE6A",x"FE69",x"FE68",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE65",x"FE65",x"FE65",
									 x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE65",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE24",x"FE25",x"FE04",x"FE05",x"FE05",
									 x"FDE4",x"FDE4",x"FDC4",x"FDC4",x"FDA4",x"FD84",x"F584",x"F564",x"FD43",x"FD23",
									 x"FCE2",x"FCC2",x"F4A2",x"F462",x"EC65",x"E4C9",x"D54E",x"D5B3",x"CDF6",x"CE17",
									 x"CE79",x"DEFB",x"E75D",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBD",
									 x"FF5B",x"FE96",x"F56E",x"EC88",x"EC25",x"F424",x"F423",x"F483",x"F4A3",x"F4C3",
									 x"FD04",x"F504",x"F524",x"FD24",x"FD44",x"FD65",x"FD65",x"FD85",x"FD85",x"FDA5",
									 x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDE5",x"FDE5",x"FE05",x"FE06",x"FE27",x"FE49",
									 x"FE4B",x"FE6C",x"FE8D",x"FEAE",x"FECF",x"FECF",x"FECF",x"FECF",x"FECF",x"FECF",
									 x"FEAF",x"FEAF",x"FEAE",x"FEAE",x"FEAE",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",
									 x"FEAC",x"FE8C",x"FE8C",x"FE8C",x"FE8B",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",
									 x"FE8A",x"FE8A",x"FE6A",x"FE69",x"FE68",x"FE68",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",x"FE45",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE65",x"FE65",x"FE65",x"FE65",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDE4",x"FDC4",x"FDC4",x"FDA4",
									 x"FDA4",x"FD84",x"FD64",x"F544",x"FD23",x"FCE3",x"FCC3",x"F4A3",x"F483",x"EC85",
									 x"E4CA",x"D52E",x"CDB3",x"C5F7",x"C619",x"CE59",x"DEDB",x"E75D",x"EF9E",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFDF",x"FFFE",x"FFFE",x"FFFE",x"FFDE",x"FF9C",x"FEB6",x"ED8F",
									 x"E4CA",x"EC46",x"F403",x"F443",x"F463",x"F483",x"FCC4",x"FCE3",x"FCE4",x"FD24",
									 x"FD24",x"FD44",x"FD65",x"FD65",x"FD85",x"FD85",x"FDA5",x"FDA6",x"FDC5",x"FDC5",
									 x"FDE5",x"FDE5",x"FDE5",x"FDE6",x"FDE6",x"FE07",x"FE08",x"FE28",x"FE29",x"FE4A",
									 x"FE6B",x"FE8C",x"FE8C",x"FEAD",x"FEAE",x"FEAE",x"FEAF",x"FEAF",x"FEAE",x"FEAE",
									 x"FEAE",x"FEAD",x"FEAD",x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",
									 x"FE8C",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE69",x"FE68",
									 x"FE68",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE25",x"FE25",x"FE45",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE25",x"FE25",x"FE25",x"FE25",x"FE05",x"FE05",x"FE05",x"FDE5",
									 x"FDE5",x"FDC5",x"FDC4",x"FDA4",x"FD84",x"FD84",x"FD64",x"FD44",x"FD44",x"FD03",
									 x"FCE3",x"FCA3",x"F483",x"EC64",x"E486",x"E4EB",x"D54F",x"CDB3",x"C616",x"C638",
									 x"CE7A",x"D6DB",x"EF5D",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFE",x"FFFF",x"FFFF",x"FFDE",x"FF7B",x"F696",x"F5F1",x"F4EA",x"F425",x"F403",
									 x"F423",x"F443",x"F483",x"FCA3",x"FCC3",x"F504",x"FD04",x"FD24",x"FD45",x"FD65",
									 x"FD65",x"FD85",x"FD85",x"FD86",x"FDA6",x"FDC5",x"FDE5",x"FDE5",x"FDE6",x"FDE7",
									 x"FDC6",x"FDE6",x"FE05",x"FE05",x"FE06",x"FE27",x"FE48",x"FE49",x"FE49",x"FE6A",
									 x"FE8B",x"FE8C",x"FEAD",x"FEAD",x"FEAD",x"FEAE",x"FEAE",x"FEAD",x"FEAD",x"FEAD",
									 x"FEAD",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FEAC",x"FE8C",x"FE8B",x"FE8B",x"FE8A",
									 x"FE8A",x"FE8A",x"FE8A",x"FE68",x"FE68",x"FE68",x"FE67",x"FE67",x"FE67",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",
									 x"FE45",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDC5",x"FDC5",x"FDA4",x"FDA4",x"FD84",
									 x"FD84",x"F564",x"F544",x"F523",x"FD03",x"F4C2",x"F482",x"F463",x"F464",x"EC66",
									 x"E4CA",x"D570",x"CDB4",x"C5F6",x"C658",x"D699",x"DEDB",x"EF5D",x"F7BE",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",
									 x"FFBD",x"FF5A",x"F6D6",x"F5D1",x"ECAA",x"EC26",x"EC23",x"F422",x"FC62",x"F483",
									 x"F4A4",x"F4C4",x"F504",x"F524",x"F525",x"FD44",x"FD43",x"FD65",x"FD85",x"FD85",
									 x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDC6",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FDE6",
									 x"FE06",x"FE06",x"FE27",x"FE27",x"FE27",x"FE48",x"FE49",x"FE69",x"FE6A",x"FE8B",
									 x"FE8B",x"FE8B",x"FE8C",x"FE8C",x"FE8C",x"FE8C",x"FE8C",x"FE8D",x"FE8C",x"FE8C",
									 x"FE8C",x"FE8B",x"FE8B",x"FE8A",x"FE8A",x"FE8A",x"FE89",x"FE89",x"FE88",x"FE68",
									 x"FE67",x"FE67",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE24",x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE05",x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDC5",
									 x"FDC4",x"FDA4",x"FDA4",x"FDA4",x"FD64",x"FD64",x"F544",x"F543",x"F503",x"FCE3",
									 x"FCC3",x"FC82",x"F483",x"EC85",x"EC87",x"E4CA",x"D54E",x"CDD4",x"CDF6",x"C637",
									 x"D699",x"DEFB",x"EF5C",x"F79E",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"FF9C",x"FF18",
									 x"F5F2",x"ED0C",x"EC87",x"F424",x"F422",x"F442",x"F483",x"F4A3",x"F4C3",x"F4E4",
									 x"F504",x"FD24",x"FD43",x"FD44",x"FD65",x"FD65",x"FD85",x"FDA5",x"FDA5",x"FDC5",
									 x"FDC5",x"FDC5",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE26",x"FE27",x"FE47",x"FE27",x"FE48",x"FE48",x"FE48",x"FE49",x"FE49",
									 x"FE6A",x"FE6A",x"FE6A",x"FE6A",x"FE6A",x"FE6A",x"FE6A",x"FE89",x"FE69",x"FE69",
									 x"FE69",x"FE69",x"FE68",x"FE68",x"FE67",x"FE67",x"FE67",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE25",x"FE25",x"FE25",x"FE24",
									 x"FE24",x"FE24",x"FE25",x"FE25",x"FE25",x"FE05",x"FE05",x"FE05",x"FE04",x"FE04",
									 x"FE04",x"FDE4",x"FDE4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FD84",x"FD84",
									 x"FD64",x"F544",x"F524",x"F504",x"F4E3",x"F4C3",x"FC83",x"F463",x"E485",x"E4A8",
									 x"DD0C",x"DD90",x"CDD4",x"D637",x"CE59",x"D69A",x"E71C",x"EF7E",x"FFBE",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FEF9",x"F613",x"F54E",x"F488",
									 x"F424",x"F422",x"F442",x"F462",x"F482",x"F4A3",x"F4C4",x"FD04",x"FD23",x"FD24",
									 x"FD44",x"FD45",x"FD64",x"FD85",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDC6",x"FDE6",
									 x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE27",x"FE27",x"FE47",x"FE48",x"FE48",x"FE48",
									 x"FE48",x"FE48",x"FE68",x"FE48",x"FE48",x"FE68",x"FE68",x"FE48",x"FE67",x"FE67",
									 x"FE67",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",x"FE45",
									 x"FE45",x"FE45",x"FE24",x"FE24",x"FE24",x"FE24",x"FE24",x"FE24",x"FE25",x"FE25",
									 x"FE05",x"FE05",x"FE05",x"FE05",x"FE04",x"FDE4",x"FDE4",x"FDC4",x"FDC4",x"FDC4",
									 x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD64",x"FD44",x"F543",x"F523",x"F503",x"F4E3",
									 x"F4A3",x"F484",x"F464",x"EC65",x"DCC8",x"DD2D",x"D592",x"CE16",x"C637",x"D679",
									 x"D6BB",x"E71D",x"EF7E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"F7FF",x"FFDF",x"FF9D",x"FEF9",x"FE34",x"F52E",x"F468",x"F424",x"F402",x"F422",
									 x"FC62",x"FC83",x"F4A3",x"FCC3",x"FCE3",x"FD24",x"FD24",x"FD44",x"FD44",x"FD64",
									 x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC6",x"FDC6",x"FDC5",x"FDC6",x"FDE6",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE26",x"FE06",
									 x"FE07",x"FE27",x"FE27",x"FE27",x"FE48",x"FE27",x"FE47",x"FE27",x"FE48",x"FE48",
									 x"FE28",x"FE48",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE24",x"FE24",x"FE24",x"FE04",x"FE04",
									 x"FE24",x"FE04",x"FE04",x"FE04",x"FE25",x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDE5",
									 x"FDE4",x"FDE4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD64",x"FD44",
									 x"FD44",x"FD23",x"FD03",x"FD02",x"FCC2",x"FCA3",x"F463",x"F444",x"EC46",x"E488",
									 x"DD2D",x"DDB2",x"D616",x"C638",x"C699",x"D6DA",x"E73C",x"EF7D",x"F7BE",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FF9D",
									 x"FF3A",x"FE96",x"F5AF",x"F4CA",x"EC46",x"EC23",x"EC22",x"F442",x"F463",x"F4A3",
									 x"F4C3",x"FCE4",x"FD04",x"FD04",x"FD24",x"FD44",x"FD64",x"FD84",x"FD84",x"FDA5",
									 x"FDA5",x"FDA5",x"FDA6",x"FDA5",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE7",
									 x"FDE7",x"FDE7",x"FDE6",x"FE06",x"FE07",x"FE07",x"FE07",x"FE07",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE28",x"FE28",x"FE28",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE24",x"FE04",x"FE04",x"FE04",x"FE04",x"FE04",x"FE04",x"FE04",
									 x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",
									 x"FD84",x"FD84",x"FD84",x"FD64",x"FD43",x"FD23",x"FD03",x"FCE3",x"FCE2",x"FCA2",
									 x"FC82",x"F463",x"EC45",x"E487",x"E4EB",x"DD4F",x"D5B3",x"CDF6",x"CE38",x"CE79",
									 x"D6FA",x"E75C",x"F79D",x"FFDE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F7DF",x"FFFF",x"FFBD",x"FEF8",x"FDF2",
									 x"F50D",x"EC66",x"EC23",x"EC22",x"F443",x"F463",x"F482",x"F4A3",x"FCC3",x"FCE3",
									 x"F503",x"FD24",x"FD44",x"F564",x"FD64",x"FD84",x"FD85",x"FD85",x"FDA5",x"FDA5",
									 x"FDA5",x"FDC5",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",
									 x"FE06",x"FE06",x"FE06",x"FE26",x"FE26",x"FE26",x"FE26",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE47",x"FE27",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE04",
									 x"FE04",x"FE04",x"FE04",x"FDE4",x"FDE4",x"FDE4",x"FDE5",x"FDE5",x"FDE4",x"FDC4",
									 x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD64",x"FD64",x"FD64",
									 x"FD23",x"FD23",x"FD03",x"FCE3",x"F4A3",x"F482",x"F463",x"F485",x"E4A8",x"DCEB",
									 x"D591",x"CDF6",x"C658",x"C67A",x"D69A",x"DEFB",x"EF5C",x"F7BE",x"FFDE",x"FFDF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"F7FF",x"F7DE",x"FF9C",x"FEF9",x"F635",x"ED4D",x"ECA8",x"F445",
									 x"F423",x"EC42",x"EC82",x"F483",x"FCC3",x"FCC3",x"FCE3",x"FD04",x"FD23",x"FD24",
									 x"FD44",x"FD44",x"FD64",x"FD85",x"FD85",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",
									 x"FDA5",x"FDC5",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE26",x"FE26",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE05",x"FE05",x"FE04",x"FE05",x"FE05",x"FDE5",x"FDE4",
									 x"FDE4",x"FDE4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FD84",x"FD83",
									 x"FD83",x"FD84",x"FD63",x"FD44",x"FD23",x"FD24",x"F504",x"F4E3",x"FCC2",x"F4A2",
									 x"F462",x"EC43",x"EC66",x"E4CA",x"DD2E",x"D592",x"CDF6",x"C638",x"C679",x"D6BB",
									 x"DF1C",x"EF5C",x"F79E",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FF9D",x"FF3B",x"F675",x"F590",x"F4EB",x"EC67",x"EC44",x"EC43",x"F443",
									 x"F482",x"F4A2",x"F4A3",x"F4C4",x"F4E3",x"F504",x"FD04",x"FD24",x"FD44",x"FD64",
									 x"FD84",x"FD65",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC6",
									 x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE26",
									 x"FE26",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE47",x"FE47",
									 x"FE47",x"FE27",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",x"FE25",
									 x"FE25",x"FE25",x"FE25",x"FE25",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FDE4",x"FDE5",x"FDE4",x"FDE4",x"FDC4",x"FDC4",x"FDE4",x"FDC4",x"FDC4",
									 x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FD64",x"FD64",x"FD44",x"FD44",x"FD24",x"FD24",
									 x"FD03",x"FD04",x"F4C3",x"F4C3",x"F4A3",x"EC84",x"EC85",x"E4A7",x"DCEC",x"D570",
									 x"CDD3",x"CE16",x"CE58",x"CE79",x"D6BA",x"E73C",x"EF7D",x"F7BE",x"FFDF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFBE",x"FF5C",
									 x"FED9",x"FE55",x"F54E",x"EC88",x"EC25",x"EC23",x"EC42",x"F462",x"F463",x"F4A3",
									 x"F4C3",x"F4C3",x"FCE4",x"FD04",x"FD24",x"FD24",x"FD44",x"FD64",x"FD64",x"FD85",
									 x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC6",x"FDC6",x"FDE6",x"FDE6",
									 x"FDE6",x"FE06",x"FDE6",x"FE06",x"FE06",x"FE06",x"FE06",x"FE27",x"FE26",x"FE26",
									 x"FE26",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE25",x"FE25",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDE4",x"FDE5",x"FDE4",
									 x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD84",x"FD84",
									 x"FD64",x"FD64",x"FD44",x"FD24",x"FD03",x"FD03",x"FCE3",x"FCC3",x"FC83",x"F462",
									 x"EC83",x"E4A6",x"E4C9",x"DD2E",x"DDD3",x"CE36",x"CE58",x"CE59",x"D6BA",x"DEFB",
									 x"EF5D",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",x"F79D",x"FF1A",x"FE55",x"F56E",
									 x"F4EA",x"EC66",x"EC23",x"EC22",x"F422",x"FC63",x"FC82",x"F4A3",x"F4C3",x"FCE3",
									 x"FD04",x"FD04",x"FD24",x"FD44",x"FD64",x"FD64",x"FD85",x"FD85",x"F585",x"FD85",
									 x"FDA5",x"FDA5",x"FDA5",x"FDC6",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE47",x"FE47",x"FE47",
									 x"FE47",x"FE47",x"FE47",x"FE47",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE47",
									 x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",
									 x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",
									 x"FDE5",x"FDE5",x"FDE4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",
									 x"FDA4",x"FD84",x"FD84",x"FD64",x"FD64",x"FD64",x"FD44",x"FD23",x"FD23",x"FD03",
									 x"FCE2",x"FCC2",x"F4A2",x"FC83",x"F463",x"F464",x"ECA7",x"E50B",x"DD4F",x"DDB3",
									 x"D617",x"CE59",x"CE99",x"D69A",x"E71C",x"EF5D",x"F79E",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFBD",x"FF5A",x"FE96",x"F5F2",x"ED2D",x"E488",x"EC45",
									 x"EC24",x"F443",x"F462",x"F463",x"F483",x"F4A3",x"FCC3",x"FCE3",x"FD04",x"FD24",
									 x"FD44",x"FD44",x"FD44",x"FD64",x"FD65",x"FD85",x"FD85",x"FD85",x"FDA5",x"FDA5",
									 x"FDA5",x"FDC5",x"FDC6",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE26",x"FE06",
									 x"FE06",x"FE26",x"FE27",x"FE27",x"FE47",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE26",x"FE26",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",
									 x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",
									 x"FDE4",x"FDE5",x"FDE5",x"FDE5",x"FDE4",x"FDE4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",
									 x"FDC4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD64",x"FD64",x"FD44",
									 x"FD44",x"FD44",x"FD23",x"FD02",x"FD03",x"FCE3",x"F4A2",x"F4A2",x"EC82",x"EC64",
									 x"EC67",x"E4C9",x"DD0D",x"DD91",x"DDF4",x"D637",x"CE59",x"CE9A",x"DEFA",x"E71B",
									 x"F77D",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDE",x"FF9D",x"F73B",x"F697",x"EDD0",x"ED2B",x"EC87",x"EC24",x"EC23",x"F442",
									 x"F462",x"F483",x"F4A3",x"FCC3",x"FCC3",x"FCE3",x"FD04",x"FD04",x"FD24",x"FD24",
									 x"FD44",x"FD64",x"FD64",x"FD65",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",
									 x"FDC5",x"FDC5",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE26",x"FE27",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE27",x"FE26",x"FE26",x"FE26",
									 x"FE27",x"FE27",x"FE27",x"FE27",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE05",x"FE05",
									 x"FE05",x"FDE5",x"FE05",x"FE05",x"FE05",x"FE05",x"FE05",x"FDE5",x"FDE5",x"FDE5",
									 x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",
									 x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD84",
									 x"FD84",x"FD63",x"FD43",x"FD43",x"FD43",x"FD23",x"FD23",x"FD03",x"FD03",x"FCC3",
									 x"FCC3",x"F484",x"F463",x"EC64",x"E484",x"E4A8",x"E50D",x"DD91",x"D5F5",x"D617",
									 x"CE59",x"D69A",x"DEDB",x"E73C",x"EF9C",x"EFBE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"FF7D",
									 x"F719",x"F695",x"F5D0",x"F50B",x"EC67",x"EC44",x"F443",x"F442",x"F463",x"F483",
									 x"F483",x"FCA3",x"FCC3",x"FCE3",x"FCE3",x"F503",x"FD03",x"FD24",x"FD24",x"FD44",
									 x"FD64",x"FD65",x"FD85",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDC5",
									 x"FDC5",x"FDC5",x"FDE5",x"FDE6",x"FDE5",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE26",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE26",x"FE27",x"FE27",x"FE27",
									 x"FE27",x"FE26",x"FE26",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE05",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",
									 x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",
									 x"FDE4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDA4",x"FDA4",x"FD84",
									 x"FD84",x"FD84",x"FD84",x"FD64",x"FD64",x"FD64",x"FD43",x"FD43",x"FD23",x"FD23",
									 x"FD03",x"F503",x"F4E3",x"FCE3",x"FCA3",x"F483",x"F484",x"F464",x"EC86",x"E4C9",
									 x"E50C",x"E56F",x"DDF3",x"D636",x"D679",x"DE9A",x"D6BB",x"DF1C",x"EF5D",x"F7BE",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"F7BD",x"F77B",x"F6D8",x"F613",
									 x"ED2D",x"EC68",x"EC45",x"EC22",x"F402",x"F422",x"F462",x"FC83",x"FC83",x"FCA3",
									 x"FCC3",x"F4E3",x"F4E3",x"FD04",x"FD04",x"FD44",x"FD44",x"FD64",x"FD65",x"FD85",
									 x"FD85",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDC5",x"FDE5",x"FDE5",
									 x"FDE5",x"FDE5",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE07",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FDE6",x"FE06",x"FDE6",
									 x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE5",x"FDE4",x"FDE4",x"FDE5",x"FDE4",x"FDC4",
									 x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",
									 x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD84",x"FD64",x"FD44",
									 x"FD44",x"FD23",x"FD23",x"FD23",x"FCE3",x"FCE3",x"FCE3",x"F4C3",x"F4A2",x"FCA2",
									 x"FC82",x"F463",x"EC64",x"EC66",x"E4CA",x"DD2E",x"DDB2",x"DE15",x"D657",x"CE79",
									 x"CE9A",x"DEDB",x"E73C",x"EF7D",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"F7DE",x"F77D",x"F6FA",x"EE55",x"F5B0",x"ED4C",x"EC87",
									 x"EC25",x"F403",x"F422",x"F442",x"F442",x"FC83",x"FC83",x"F4A3",x"F4C4",x"F4E4",
									 x"F4E3",x"F503",x"F523",x"FD44",x"FD44",x"FD64",x"FD64",x"FD64",x"FD84",x"FD84",
									 x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDA5",x"FDC5",x"FDC5",x"FDC5",x"FDE6",
									 x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",
									 x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FE06",x"FDE6",
									 x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE5",x"FDE5",x"FDC5",x"FDE5",x"FDE5",x"FDE5",
									 x"FDC5",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDC4",x"FDA4",x"FDC4",x"FDC4",x"FDA4",
									 x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FD83",x"FD84",
									 x"FD84",x"FD64",x"FD64",x"FD64",x"F563",x"F543",x"FD23",x"FD03",x"FD03",x"FCE3",
									 x"FCC4",x"FCC4",x"FCA3",x"FC83",x"F462",x"F462",x"EC63",x"EC85",x"E4C8",x"DCEB",
									 x"E570",x"DDD5",x"D616",x"D678",x"D6BA",x"D6DC",x"DF1D",x"E75E",x"EF9E",x"FFDF",
									 x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",x"F7DE",
									 x"F7BF",x"FFBE",x"FF7C",x"F719",x"F6B6",x"EDB0",x"ECEC",x"EC89",x"EC65",x"F443",
									 x"F423",x"F443",x"FC63",x"F483",x"F4A3",x"F4A3",x"F4C3",x"F4C3",x"F4E3",x"F503",
									 x"F524",x"FD24",x"FD44",x"FD44",x"FD44",x"FD44",x"FD64",x"FD85",x"FD85",x"FD85",
									 x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC6",x"FDC6",
									 x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",
									 x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",
									 x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE5",x"FDE5",x"FDC5",x"FDC5",x"FDC5",
									 x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC4",x"FDA4",x"FDA4",x"FDA4",
									 x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FDA4",x"FD84",
									 x"FD84",x"FD84",x"FD84",x"FD64",x"FD63",x"FD63",x"FD63",x"FD63",x"FD43",x"F543",
									 x"F523",x"F523",x"F503",x"F4E3",x"FCC3",x"FCA3",x"F4A2",x"F482",x"F483",x"F484",
									 x"EC45",x"E466",x"DCA9",x"DD2D",x"DD91",x"DDF3",x"DE56",x"D699",x"D699",x"D6BA",
									 x"DEFB",x"E75D",x"F79E",x"F7BF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFE",x"FFFE",x"FFFF",x"FFDF",x"FFBE",x"F7BE",
									 x"FF9C",x"FF1A",x"F656",x"F5F2",x"ED4D",x"ECA8",x"E446",x"EC24",x"F423",x"F442",
									 x"F442",x"F463",x"F483",x"F4A3",x"F4C3",x"F4E3",x"FCE4",x"FD03",x"FD03",x"FD04",
									 x"FD24",x"FD24",x"FD44",x"FD64",x"FD64",x"FD65",x"FD65",x"FD65",x"FD85",x"FD84",
									 x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA6",x"FDA5",x"FDC6",x"FDC6",x"FDA5",x"FDC5",
									 x"FDC5",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",
									 x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDE6",x"FDE6",x"FDE6",x"FDE6",x"FDE5",x"FDC5",
									 x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",
									 x"FDA5",x"FDA5",x"FDA5",x"FDA4",x"FDA4",x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",
									 x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",x"FD64",x"FD64",x"FD64",x"FD44",x"FD44",
									 x"FD43",x"FD43",x"FD23",x"FD23",x"F503",x"F503",x"F4E2",x"F4E2",x"F4C2",x"F4A3",
									 x"F483",x"F483",x"EC82",x"EC62",x"E463",x"E486",x"E4CA",x"E52E",x"DD92",x"DE16",
									 x"D658",x"D658",x"D699",x"D6DA",x"DEFB",x"EF5C",x"F79D",x"FFBE",x"FFBF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDE",x"F7DE",x"FFDE",x"FF9D",x"FF1B",x"FEB8",
									 x"EE33",x"ED4E",x"ECCB",x"EC68",x"EC05",x"F403",x"F422",x"F422",x"F442",x"F462",
									 x"F482",x"F4A3",x"F4A3",x"F4C3",x"F4E4",x"FCE4",x"FD04",x"FD04",x"FD24",x"FD44",
									 x"FD44",x"FD44",x"FD45",x"FD65",x"FD65",x"FD64",x"FD84",x"FD85",x"FD85",x"FD85",
									 x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",
									 x"FDC5",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC6",x"FDC5",x"FDC5",x"FDC6",
									 x"FDC6",x"FDC6",x"FDC6",x"FDE6",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDC5",x"FDA5",
									 x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA4",x"FDA4",x"FDA4",x"FD84",
									 x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",x"FD64",x"FD64",x"FD64",
									 x"FD64",x"FD44",x"FD43",x"FD43",x"FD23",x"FD23",x"FD03",x"FD04",x"FD04",x"FCE4",
									 x"FCE4",x"F4C3",x"FCC3",x"FCC2",x"FC82",x"F462",x"F462",x"F443",x"EC65",x"EC66",
									 x"E487",x"E4EB",x"DD6F",x"D5D3",x"DE35",x"D678",x"D69A",x"D69A",x"DEBA",x"E6DB",
									 x"E73C",x"EF9D",x"FFBE",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDF",x"FFDF",x"FFDE",x"FFDE",x"FFBE",x"FF9D",x"FF7C",x"FEF8",x"F676",x"F5B2",
									 x"ED0D",x"EC88",x"EC46",x"EC24",x"EC24",x"EC23",x"F443",x"F463",x"F483",x"F483",
									 x"F4A3",x"F4A3",x"F4C3",x"F4E3",x"F504",x"FD04",x"FD04",x"F504",x"FD25",x"FD25",
									 x"FD24",x"FD44",x"FD64",x"FD64",x"FD64",x"FD65",x"FD65",x"FD65",x"FD85",x"FD85",
									 x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC5",
									 x"FDC5",x"FDC5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDC5",x"FDC5",x"FDA5",x"FDA5",
									 x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FD85",x"FD85",
									 x"FD85",x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",x"FD64",x"FD64",x"FD64",
									 x"FD64",x"FD64",x"FD64",x"F564",x"F564",x"F544",x"FD44",x"FD23",x"FD23",x"FD23",
									 x"FD03",x"FD03",x"FCE3",x"FCE4",x"F4C4",x"F4C3",x"F4A3",x"F482",x"F482",x"F483",
									 x"F463",x"EC44",x"EC45",x"EC66",x"E4AA",x"E50D",x"E570",x"E5F3",x"E697",x"DE78",
									 x"D678",x"DEBA",x"DEFB",x"E71C",x"EF5D",x"FFBE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDF",x"FFDF",x"FFDF",x"FFBE",x"F77C",x"F71A",x"F676",x"F5F2",x"F58E",x"ED0B",
									 x"EC88",x"EC66",x"F444",x"F423",x"F422",x"F463",x"F463",x"F463",x"F483",x"F4A3",
									 x"F4C3",x"F4C3",x"F4E3",x"F4E4",x"F504",x"F504",x"FD04",x"FD23",x"FD24",x"FD44",
									 x"FD44",x"FD44",x"FD45",x"FD44",x"FD65",x"FD65",x"FD65",x"FD65",x"FD85",x"FD85",
									 x"FD85",x"FD85",x"FD85",x"FD85",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FD85",x"FDA5",
									 x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FDA5",x"FD85",x"FD84",x"FD84",
									 x"FD84",x"FD84",x"FD84",x"FD84",x"FD84",x"FD64",x"FD64",x"FD64",x"FD64",x"FD64",
									 x"FD64",x"FD64",x"FD64",x"FD44",x"FD44",x"FD44",x"FD43",x"FD43",x"FD43",x"F544",
									 x"F544",x"F523",x"F523",x"F503",x"F503",x"F503",x"F4E2",x"F4C2",x"F4A3",x"F4A3",
									 x"F483",x"F483",x"F463",x"EC43",x"F463",x"F464",x"EC86",x"E4C9",x"E4EB",x"E52D",
									 x"DDB2",x"DDF4",x"D636",x"D678",x"DEDB",x"DEFC",x"DF1C",x"E73C",x"EF5D",x"F79D",
									 x"F7BE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"F7DF",
									 x"F7DF",x"F79E",x"FF5C",x"F719",x"F6B7",x"EDD2",x"E52E",x"ECCA",x"EC67",x"EC24",
									 x"F403",x"EC43",x"F443",x"F443",x"F443",x"F463",x"F483",x"F4A2",x"F4C2",x"F4E3",
									 x"F503",x"F503",x"F503",x"F503",x"F503",x"F524",x"F524",x"F524",x"F524",x"FD24",
									 x"FD44",x"FD44",x"FD44",x"FD45",x"FD65",x"FD65",x"FD65",x"FD85",x"FD85",x"FD84",
									 x"FD85",x"FD85",x"FD85",x"FD85",x"FD84",x"FD64",x"FD64",x"FD65",x"FD85",x"FD85",
									 x"FD85",x"FD65",x"FD85",x"FD65",x"FD64",x"FD64",x"FD64",x"FD64",x"FD64",x"FD64",
									 x"FD64",x"FD64",x"FD64",x"FD64",x"FD64",x"FD43",x"F543",x"F543",x"F543",x"F523",
									 x"FD24",x"FD24",x"FD23",x"FD23",x"FD03",x"FD03",x"FCE3",x"FCE3",x"F503",x"F4E2",
									 x"F4E3",x"F4E2",x"F4C2",x"F4A2",x"F482",x"F462",x"F462",x"F463",x"EC64",x"E465",
									 x"EC46",x"E488",x"E4CB",x"DD4F",x"D5B2",x"D635",x"D677",x"D699",x"D699",x"D6BA",
									 x"D6FB",x"DF3D",x"EF5D",x"F79E",x"F7BE",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"F7DF",x"F7BF",x"F77D",
									 x"F75C",x"F6FA",x"F698",x"F634",x"ED90",x"ED0C",x"ECCA",x"EC67",x"EC46",x"F425",
									 x"F424",x"F423",x"F443",x"F462",x"F483",x"F482",x"F482",x"F4A3",x"F4C3",x"F4C3",
									 x"F4C3",x"F4E4",x"F504",x"F504",x"F504",x"FD24",x"FD24",x"FD24",x"FD24",x"FD44",
									 x"FD44",x"FD45",x"FD45",x"FD65",x"FD44",x"FD44",x"FD64",x"FD64",x"FD44",x"FD44",
									 x"FD44",x"FD44",x"FD64",x"FD64",x"FD65",x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",
									 x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",x"FD44",x"FD43",x"FD43",x"FD43",
									 x"FD23",x"F523",x"F523",x"F523",x"F503",x"F503",x"F503",x"F503",x"FCE3",x"FCE3",
									 x"FCE3",x"FCC3",x"FCC3",x"FCA3",x"F4A3",x"F4A3",x"F4A3",x"F4A3",x"F483",x"EC63",
									 x"EC63",x"F463",x"F444",x"EC45",x"EC88",x"E4EB",x"DD0E",x"DD70",x"E5D3",x"DE36",
									 x"D657",x"CE98",x"D6DA",x"D6FB",x"DF1B",x"E73C",x"EF5D",x"EF7D",x"F7BE",x"FFDF",
									 x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"F7DF",x"FFDF",x"FFDF",x"FF9E",x"FF7C",
									 x"FF1A",x"F676",x"EE14",x"F5B0",x"F52D",x"ECCB",x"EC89",x"EC67",x"EC45",x"EC45",
									 x"EC44",x"F423",x"F443",x"F443",x"F463",x"F463",x"F483",x"F483",x"F4A3",x"F4C3",
									 x"F4C3",x"F4C3",x"FCE3",x"FCE3",x"FCE4",x"F504",x"F504",x"FD04",x"FD04",x"FD04",
									 x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",
									 x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD24",x"FD04",x"FD04",x"FD24",x"FD24",
									 x"FD24",x"FD24",x"FD23",x"FD03",x"FD03",x"FD03",x"FD03",x"F503",x"F503",x"F4E3",
									 x"F4E3",x"F4E3",x"F4C3",x"F4C3",x"F4A3",x"F4A3",x"F4A3",x"F4A3",x"F483",x"F463",
									 x"F463",x"F464",x"F444",x"EC65",x"EC66",x"EC66",x"E486",x"E4A8",x"E4EA",x"E52D",
									 x"E570",x"E5D2",x"DE56",x"DE78",x"E6DA",x"E6DB",x"E6FB",x"E71B",x"E73C",x"E75C",
									 x"EF7D",x"FFBE",x"FFDF",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFDF",x"FFDF",x"FFBE",x"F7BE",x"F7BE",x"EF7D",x"EF5C",x"F75C",x"F71A",
									 x"F6B8",x"F635",x"F5D1",x"F54D",x"E4EA",x"ECA9",x"EC67",x"EC25",x"F424",x"F423",
									 x"F423",x"F443",x"F463",x"FC63",x"F463",x"F483",x"F483",x"F483",x"F4A3",x"F4A3",
									 x"F4C3",x"F4C3",x"F4C3",x"FCE4",x"FCE4",x"FCE4",x"FCE4",x"F504",x"FD03",x"FD04",
									 x"FD04",x"FD04",x"FD04",x"FD04",x"FD04",x"FD04",x"FD04",x"FD04",x"F504",x"FD04",
									 x"FD04",x"FD04",x"FD04",x"FD04",x"FD04",x"FD04",x"FD04",x"FD04",x"FCE3",x"FCE3",
									 x"FCE3",x"FCE3",x"FCE3",x"F4C3",x"F4C3",x"F4C3",x"F4A3",x"F4A3",x"F483",x"F483",
									 x"F483",x"F483",x"F483",x"F463",x"EC63",x"EC63",x"F444",x"EC45",x"EC66",x"E487",
									 x"E4A9",x"E4EA",x"E52D",x"E590",x"DE14",x"DE57",x"DE79",x"DE99",x"DEB8",x"DEBA",
									 x"E6FB",x"E71D",x"E73D",x"EF7D",x"F7BE",x"F7BE",x"FFBF",x"FFDF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDE",
									 x"FFDF",x"FFFF",x"FFFF",x"F7DF",x"F7DE",x"F79E",x"F75C",x"F6FA",x"F6B8",x"F675",
									 x"EE13",x"F5D1",x"ED6F",x"ED0C",x"ECC9",x"EC87",x"EC66",x"EC45",x"EC44",x"F444",
									 x"F443",x"F442",x"F442",x"F442",x"F443",x"F463",x"F483",x"F483",x"F4A3",x"F4A3",
									 x"F4A3",x"F4C3",x"F4C3",x"F4C3",x"F4C3",x"F4C3",x"F4C3",x"F4E3",x"F4E3",x"F4E3",
									 x"F4E3",x"F4E3",x"F4E4",x"F4E4",x"F4C4",x"F4E4",x"F4E4",x"F4E3",x"F4E3",x"F4E3",
									 x"F4E3",x"F4E3",x"F4C3",x"F4C3",x"FCC3",x"F4C3",x"F4A3",x"F4A3",x"F4A3",x"F483",
									 x"F483",x"F482",x"F482",x"F463",x"F462",x"F462",x"F462",x"F463",x"EC64",x"EC64",
									 x"EC85",x"ECA6",x"ECA8",x"ECC9",x"E4EB",x"E54D",x"E590",x"E5D2",x"DDF4",x"DE36",
									 x"DE78",x"D6BB",x"DEFC",x"DF1C",x"E71B",x"E73C",x"EF5D",x"EF7E",x"EF7E",x"F7BE",
									 x"F7BE",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F7DF",
									 x"F7DF",x"FFDE",x"FFBE",x"F79D",x"FF9D",x"FF7C",x"F75C",x"FF3A",x"F6D8",x"F655",
									 x"F5F2",x"ED6F",x"ED2D",x"E4EA",x"E4A9",x"E488",x"E466",x"EC45",x"EC44",x"F424",
									 x"EC24",x"F424",x"F444",x"F463",x"F463",x"F463",x"F483",x"F483",x"F483",x"F483",
									 x"F483",x"F483",x"FC83",x"FC83",x"FC83",x"F4A3",x"F4A3",x"F4A3",x"FCA3",x"FCA3",
									 x"F4A3",x"F4A3",x"F4A3",x"F4A3",x"F483",x"F483",x"F483",x"FC84",x"F464",x"F484",
									 x"F483",x"F483",x"F483",x"F463",x"F463",x"F464",x"F463",x"EC43",x"EC64",x"EC44",
									 x"EC44",x"EC65",x"EC66",x"EC87",x"E4A8",x"E4AA",x"E4EC",x"E52D",x"E570",x"E5B2",
									 x"E5F4",x"E657",x"E699",x"E6DA",x"E6DA",x"E6DA",x"E6DA",x"E6FB",x"E71C",x"EF5D",
									 x"EF9D",x"F79E",x"F7BE",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"F7DF",x"F7DF",
									 x"F7DF",x"FFDF",x"FFBE",x"F7BD",x"F77C",x"F73B",x"F71A",x"F6F9",x"F6B8",x"F676",
									 x"F634",x"EDF2",x"ED90",x"ED4E",x"ED0C",x"ECEA",x"ECA9",x"ECA8",x"EC87",x"F466",
									 x"F445",x"EC64",x"EC64",x"EC44",x"EC44",x"F424",x"F424",x"F423",x"F443",x"F443",
									 x"F443",x"F443",x"F463",x"F463",x"F442",x"F462",x"F462",x"F462",x"F462",x"F442",
									 x"F443",x"F443",x"F443",x"F443",x"F444",x"F444",x"F443",x"F443",x"EC44",x"EC44",
									 x"EC66",x"EC66",x"F466",x"EC87",x"ECA8",x"E4C9",x"E4EA",x"E52B",x"E54E",x"E58F",
									 x"E5B1",x"EDF3",x"EE55",x"EE56",x"E678",x"E698",x"DE99",x"E6DB",x"E6FC",x"E71D",
									 x"EF3C",x"EF5D",x"EF7D",x"EF7D",x"F79E",x"F7BE",x"F7DF",x"FFDF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"F7BF",x"F7DE",
									 x"F7BE",x"F7BE",x"F7BE",x"F79E",x"EF7D",x"F75C",x"EF1A",x"EEB8",x"E656",x"EE35",
									 x"EDF3",x"EDD1",x"E56F",x"E52D",x"ECEC",x"ECCB",x"ECAA",x"ECA9",x"EC88",x"EC66",
									 x"F445",x"F444",x"F423",x"F423",x"F442",x"F442",x"F422",x"F422",x"F422",x"F422",
									 x"EC22",x"F422",x"F422",x"EC22",x"F422",x"F422",x"F441",x"EC42",x"EC42",x"EC43",
									 x"EC63",x"EC64",x"EC45",x"EC45",x"EC66",x"EC67",x"EC89",x"ECAA",x"E4CB",x"E4EC",
									 x"E50E",x"DD4F",x"DD91",x"DDD2",x"D5F4",x"DE36",x"DE77",x"E6B9",x"E6FB",x"E6FB",
									 x"DF1B",x"E71B",x"E71B",x"E73B",x"E73C",x"EF7C",x"EF7D",x"EF9E",x"F7BE",x"F7BE",
									 x"FFDF",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFE",x"FFDE",x"FFDE",x"FFDE",x"FFDF",x"FFDF",x"F7DF",x"F7DF",x"F7DF",x"F7DF",
									 x"F7BF",x"F79D",x"EF7D",x"EF5C",x"EF5B",x"F75B",x"F73A",x"F6F8",x"EEB7",x"EE76",
									 x"EE14",x"EDD2",x"E571",x"ED4F",x"E52E",x"E4EC",x"E4CA",x"E4C8",x"E4A7",x"EC66",
									 x"F446",x"F426",x"F425",x"F425",x"F425",x"F424",x"EC24",x"EC04",x"EC24",x"EC04",
									 x"EC04",x"EC24",x"EC45",x"EC45",x"EC66",x"EC66",x"EC67",x"E488",x"DCA9",x"E4CA",
									 x"E4EB",x"E52D",x"E54F",x"E590",x"E5B2",x"E5F3",x"E635",x"E656",x"DE78",x"DEB8",
									 x"DED9",x"DEDA",x"DEFA",x"DF1B",x"E73C",x"E75D",x"E77E",x"EF7E",x"EF7E",x"F79E",
									 x"F79E",x"FFBF",x"F7BF",x"F7DF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"F7DF",x"FFDF",x"FFDE",x"F7BE",
									 x"F7BE",x"F7DE",x"F7DE",x"F7BD",x"F79C",x"F77C",x"F73B",x"F6FA",x"EED9",x"EED8",
									 x"EEB7",x"EE96",x"EE56",x"EE35",x"EE14",x"EDF3",x"EDF3",x"EDD2",x"EDD2",x"EDD2",
									 x"F5B2",x"EDB1",x"EDD0",x"EDD0",x"F5D0",x"EDD0",x"EDB0",x"EDD0",x"EDD1",x"EDD2",
									 x"EDD2",x"EDD3",x"EDD3",x"EDD4",x"E614",x"E634",x"E634",x"DE55",x"DE76",x"E697",
									 x"E6B8",x"E6B9",x"E6FA",x"E71B",x"E73C",x"E73C",x"EF5D",x"EF5D",x"EF5D",x"EF7D",
									 x"F79D",x"F79D",x"F7BE",x"F7DF",x"F7DF",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFDF",x"FFDF",x"FFFF",x"FFDF",x"FFDF",x"FFDF",x"F7DF",x"F7DF",x"F7DF",x"F7BE",
									 x"F7BE",x"F7BE",x"F79D",x"F79D",x"F79D",x"F79D",x"F79D",x"F79D",x"F77D",x"F77D",
									 x"F75D",x"EF5C",x"EF5C",x"EF5C",x"EF5C",x"EF5C",x"EF5C",x"EF5C",x"EF3C",x"EF3C",
									 x"EF3C",x"EF3C",x"EF3C",x"EF3C",x"EF3B",x"EF3B",x"EF3B",x"EF3C",x"EF3C",x"EF3C",
									 x"EF3B",x"E73B",x"E73B",x"E73B",x"E73B",x"E73C",x"E71B",x"E73C",x"EF5D",x"EF7D",
									 x"EF7E",x"F79E",x"F79E",x"F7BF",x"F7BF",x"FFDF",x"FFDE",x"FFDE",x"FFFE",x"FFFE",
									 x"FFFE",x"FFFE",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"F7BE",x"F7BE",
									 x"F7BE",x"F7BE",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"EF9E",x"EF7D",x"EF7D",
									 x"EF7D",x"EF7D",x"EF7D",x"EF7E",x"EF7E",x"EF7E",x"EF7E",x"EF7E",x"EF7E",x"EF5E",
									 x"EF5D",x"EF5D",x"EF5D",x"EF7D",x"EF7D",x"EF7D",x"EF5D",x"EF5D",x"EF7D",x"EF7D",
									 x"EF7D",x"F79E",x"F79E",x"F79E",x"F79E",x"F79E",x"F7BE",x"F7BE",x"FFDF",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDF",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",
									 x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F79E",x"F79E",x"F7BE",x"F7BE",x"F7BE",
									 x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"F7BE",x"FFDF",x"FFDF",x"FFDF",x"FFDF",
									 x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFDF",
									 x"FFDF",x"FFDF",x"FFDF",x"FFDF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",
									 x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"FFFF");

	------------------------------------------------------------------------------------------------
	-- Internal signals	
	------------------------------------------------------------------------------------------------	
	-- Counter
	signal cntH : integer range 0 to imSizeH_g - 1;
	signal cntV : integer range 0 to imSizeV_g - 1;

	-- Color Generation
	signal color         : std_logic_vector(15 downto 0) := "1111100000000000"; -- Start with red

begin	
	-- Strobe out can be always high, data is sent on every clock 
	strobe_out <= '1' when resetn = '1' else '0';

	-- Set the image output signals
	row_out <= to_unsigned(cntH, rowSize_g);
	col_out <= to_unsigned(cntV, colSize_g);
	d_out   <= color;
	
	------------------------------------------------------------------------------------------------
	-- Read process
	------------------------------------------------------------------------------------------------
	rom_read : process(clk)
	begin
		-- Wait till the next rising edge occures
		if (rising_edge(clk)) then
			-- Read the requested data
			color <= blockrom(cntH + cntV * imSizeH_g);
		end if;
	end process rom_read;
	
	------------------------------------------------------------------------------------------------
	-- Row and Column process
	-- This process creates the signals to loop through all pixels
	------------------------------------------------------------------------------------------------
	changeRowColumn : process(clk)
	begin
		if rising_edge(clk) then
			if (resetn = '0') then
				-- Reset everything
				cntH <= 0;
				cntV <= 0;
			else
				-- Increment the row and column			
				if (cntH = imSizeH_g - 1) then
					cntH <= 0;
					if (cntV = imSizeV_g - 1) then
						cntV <= 0;
					else
						cntV <= cntV + 1;
					end if;
				else
					cntH <= cntH + 1;
				end if;
			end if;
		end if;
	end process changeRowColumn;
end architecture RTL;
