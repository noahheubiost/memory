-- # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # #
-- #                                                                     #
-- #      Hardware description by Lukas Leuenberger l1leuenb@hsr.ch      #
-- #                                                                     #
-- #                            Created: 12.12.2019                      #
-- #                        Last modified: 12.12.2019                     #
-- #                                                                     #
-- #          Copyright by Hochschule fuer Technik in Rapperswil         #
-- #                                                                     #
-- #                                                                     #
-- # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # # #

------------------------------------------------------------------------------------------------
-- Library declarations
------------------------------------------------------------------------------------------------
-- Standard library ieee	
library ieee;
-- This package defines the basic std_logic data types and a few functions.								
use ieee.std_logic_1164.all;
-- This package provides arithmetic functions for vectors.		
use ieee.numeric_std.all;
-- This package provides functions for the calcualtion with real values.
use ieee.math_real.all;
-- This package provides file specific functions.
use std.textio.all;
-- This package provides file specific functions for the std_logic types.
use ieee.std_logic_textio.all;

------------------------------------------------------------------------------------------------
-- Entity declarations
------------------------------------------------------------------------------------------------
entity compImage is
	generic(
		imSizeH_g : integer := 256; --output picture size
		imSizeV_g : integer := 256; --output picture size
		imSizeCompTotal_g : integer := 27780; --picture rom size
		-- bus size
		rowSize_g         : integer := 8;
		colSize_g         : integer := 8
	);
	port(
		-- Reset und Clock
		resetn     : in  std_logic;     -- Synchronous Negative Reset
		clk        : in  std_logic;     -- Clock
		-- FPGA Image out
		row_out    : out unsigned(rowSize_g - 1 downto 0);
		col_out    : out unsigned(colSize_g - 1 downto 0);
		d_out      : out std_logic_vector(15 downto 0);
		strobe_out : out std_logic
	);
end entity compImage;

---------------------------------------------------------------------
-- Architecture declarations
---------------------------------------------------------------------
architecture RTL of compImage is
	------------------------------------------------------------------------------------------------
	-- internal types
	------------------------------------------------------------------------------------------------
	type rom_type is array (0 to (imSizeCompTotal_g)) of std_logic_vector(17 downto 0);

	------------------------------------------------------------------------------------------------
	-- Internal constants
	------------------------------------------------------------------------------------------------
	constant blockrom : rom_type := (x"0FFFF",x"100FE",x"20003",x"0FFFF",x"10074",x"0FFFE",x"0FFFF",x"10087",x"0FFFF",x"100FE",
									 x"0FFFF",x"1006B",x"0FFFE",x"0FFBE",x"0FFBD",x"0FF9D",x"0F79C",x"0F77C",x"0FF7C",x"0FF5B",
									 x"0FF3A",x"0FF1A",x"0FF19",x"0FEF9",x"0FEF8",x"10000",x"0FED7",x"10003",x"0FEF7",x"10001",
									 x"0FED7",x"10000",x"0FED8",x"10000",x"0FEF9",x"0FF19",x"10000",x"0FF1A",x"10000",x"0FF5B",
									 x"0F77C",x"10000",x"0FF7B",x"0FF9C",x"0FFBD",x"10000",x"0FFFE",x"0FFFF",x"1006A",x"0FFFF",
									 x"10065",x"0FFDF",x"0FFDE",x"0FFBE",x"10000",x"0FFBD",x"10000",x"0F77B",x"0F719",x"0F6D7",
									 x"0F676",x"0F613",x"0F5F2",x"0F5B0",x"0F58F",x"0F54E",x"0F52D",x"0F50C",x"0ECEB",x"0ECAA",
									 x"0ECA9",x"0EC88",x"0EC68",x"0F447",x"10004",x"0EC67",x"0EC68",x"0EC88",x"0ECA9",x"0F4AA",
									 x"0F4CA",x"0F4EB",x"0F52C",x"0F54D",x"0F58F",x"0F5B0",x"0FDD1",x"0F613",x"0F675",x"0FEB7",
									 x"0F6F9",x"0FF3A",x"0FF9C",x"0FF9D",x"0FFBE",x"10000",x"0FFDE",x"0FFFF",x"10065",x"0FFFF",
									 x"10064",x"0FFDF",x"0FFBD",x"0FF7C",x"0FF3B",x"0FF19",x"0F6D7",x"0F6B6",x"0F654",x"0F5F2",
									 x"0F5B0",x"0F56E",x"0F50C",x"0ECEC",x"0F4EB",x"0F4C9",x"0EC88",x"0EC67",x"0F446",x"0F425",
									 x"0F405",x"0F404",x"10000",x"0F403",x"0F402",x"0EBE2",x"10003",x"0F3E2",x"0F3E3",x"10000",
									 x"0F404",x"10000",x"0F424",x"0F425",x"0F467",x"0F488",x"0F4A9",x"0F4CA",x"0F4EB",x"0F50D",
									 x"0F54F",x"0F590",x"0F5D2",x"0F634",x"0FE76",x"0FEB8",x"0FEF9",x"0FF3B",x"0FF7C",x"0FFBD",
									 x"0FFFE",x"0FFFF",x"10063",x"0FFFF",x"1005D",x"0FFDF",x"10001",x"0FFDE",x"0FFBD",x"0FF9C",
									 x"0FF9B",x"0FF5A",x"0FED8",x"0FE96",x"0FE54",x"0FE12",x"0FDB0",x"0F56E",x"0F50C",x"0F4CA",
									 x"0F4A9",x"0F488",x"0EC68",x"0EC47",x"0EC46",x"0EC45",x"0EC24",x"0EC04",x"10000",x"0EBE3",
									 x"10000",x"0EC03",x"10000",x"0EBE3",x"0F3E2",x"10004",x"0EC03",x"10002",x"0EC04",x"10002",
									 x"0EC25",x"0EC26",x"0EC47",x"10000",x"0EC67",x"0F488",x"0F4A9",x"0F4CB",x"0F50C",x"0F54E",
									 x"0F5B0",x"0FDF2",x"0FE34",x"0FE75",x"0FED7",x"0FF19",x"0FF9C",x"0FFBD",x"0FFDD",x"0FFDE",
									 x"0FFFF",x"1005F",x"0FFFF",x"1005A",x"0FFFE",x"10000",x"0FFDE",x"0FFBD",x"0FF7C",x"0FF3A",
									 x"0FEF8",x"0FE96",x"0F634",x"0FDF1",x"0F56F",x"0ED2D",x"0ECEB",x"0ECCA",x"0EC88",x"0F467",
									 x"0F446",x"0F425",x"10000",x"0F424",x"10000",x"0F403",x"0F423",x"10000",x"0F422",x"0FC22",
									 x"10000",x"0F402",x"10000",x"0F422",x"0FC22",x"10000",x"0F422",x"0F442",x"10008",x"0F422",
									 x"10003",x"0F423",x"10000",x"0F403",x"0F423",x"0EC24",x"10000",x"0EC25",x"10000",x"0EC46",
									 x"0EC67",x"0EC88",x"0ECAA",x"0ECEB",x"0ED0D",x"0F56F",x"0F5F2",x"0EE34",x"0F696",x"0FEF8",
									 x"0FF5A",x"0FF9C",x"0FFBD",x"0FFDD",x"0FFDE",x"0FFFE",x"0FFFF",x"10059",x"0FFFF",x"10058",
									 x"0FFFE",x"0FFDE",x"0FFBD",x"0F75C",x"0FF3A",x"0F6D8",x"0F675",x"0F5F2",x"0F5B0",x"0F52D",
									 x"0F4CB",x"0F489",x"0EC47",x"0F446",x"0F425",x"0F424",x"0EC03",x"0EC23",x"0F403",x"0F402",
									 x"0F422",x"10000",x"0F443",x"10001",x"0F463",x"10003",x"0FC83",x"0F483",x"1000C",x"0FC83",
									 x"10000",x"0F463",x"10002",x"0F443",x"10000",x"0F462",x"10000",x"0F442",x"10000",x"0F422",
									 x"0F402",x"0F403",x"10000",x"0F424",x"0EC25",x"0EC47",x"0EC48",x"0F469",x"0F4AA",x"0F52D",
									 x"0F590",x"0FDF2",x"0FE34",x"0F6B7",x"0F719",x"0F73A",x"0F77C",x"0F7BE",x"0FFFF",x"10058",
									 x"0FFFF",x"10057",x"0FFDE",x"0FF9D",x"0FF3B",x"0FEB8",x"0FE55",x"0FDF1",x"0F56D",x"0ED0B",
									 x"0ECC9",x"0EC88",x"0EC66",x"0F445",x"0F424",x"0F403",x"0EC03",x"0EC23",x"0F423",x"0EC22",
									 x"0F422",x"10000",x"0F442",x"0F463",x"10001",x"0F482",x"0F483",x"0F4A3",x"0F483",x"0F4A3",
									 x"10002",x"0F4C3",x"1000D",x"0F4A3",x"10005",x"0F482",x"0F462",x"0F442",x"0F462",x"0F442",
									 x"10000",x"0F422",x"0EC22",x"0F422",x"0F423",x"10000",x"0F403",x"0F424",x"0F425",x"0F446",
									 x"0F467",x"0F4A9",x"0F4EB",x"0FD4E",x"0FDD1",x"0FE53",x"0FEB7",x"0FF5A",x"0FFBD",x"0FFDE",
									 x"0FFFF",x"10056",x"0FFFF",x"10054",x"0FFDE",x"0FF7C",x"0FF3A",x"0FED7",x"0FE55",x"0F5D2",
									 x"0F54E",x"0ECEC",x"0ECA9",x"0EC66",x"0E425",x"0EC24",x"10000",x"0EC03",x"10000",x"0EC22",
									 x"0F422",x"0F443",x"0F463",x"10001",x"0FC83",x"10001",x"0F4A3",x"10001",x"0F4C3",x"0FCC3",
									 x"0F4C3",x"0FCC3",x"10000",x"0FCE4",x"10001",x"0F4E4",x"10008",x"0FCE4",x"10001",x"0FCE3",
									 x"0F4E3",x"0F4C3",x"0F4E3",x"10002",x"0F4C3",x"10000",x"0FCC3",x"0F4A3",x"10000",x"0FCA3",
									 x"0FC83",x"0F483",x"10000",x"0F463",x"10001",x"0F443",x"0F422",x"10000",x"0EC02",x"0EC03",
									 x"10000",x"0EC24",x"0EC25",x"0EC67",x"0ECA9",x"0ECEB",x"0ED4E",x"0EDD1",x"0F634",x"0F696",
									 x"0FF19",x"0FF7B",x"0FFBD",x"0FFFF",x"10053",x"0FFFF",x"10050",x"0FFDF",x"0FFBE",x"0FF9D",
									 x"0FF5B",x"0FEF8",x"0F655",x"0F5F1",x"0F54D",x"0ECCA",x"0EC48",x"0EC26",x"0EC04",x"0EC03",
									 x"0EC02",x"0F402",x"0F422",x"10001",x"0F442",x"0F463",x"10000",x"0F483",x"0F4A3",x"10002",
									 x"0FCA3",x"0FCC4",x"10000",x"0FCE4",x"10004",x"0FD04",x"10011",x"0F504",x"0FD04",x"10004",
									 x"0FCE4",x"0FCC3",x"0FCC4",x"10001",x"0FCC3",x"10000",x"0FCA3",x"0F4A3",x"10000",x"0F483",
									 x"10000",x"0F462",x"10000",x"0F442",x"0F422",x"0EC22",x"10000",x"0EBE2",x"0EC03",x"0EC04",
									 x"0EC45",x"0E467",x"0ECC9",x"0F52D",x"0F5B0",x"0FE34",x"0FEB7",x"0FF5B",x"0FF9D",x"0FFBE",
									 x"0FFFE",x"0FFFF",x"0F7FF",x"0FFFF",x"1004D",x"0FFFF",x"1004F",x"0FFDF",x"0F79D",x"0FF3A",
									 x"0F6B7",x"0F633",x"0F590",x"0F50C",x"0F4A9",x"0EC67",x"0EC45",x"0F424",x"0F423",x"0F422",
									 x"10000",x"0F442",x"10000",x"0F462",x"10000",x"0F463",x"0F483",x"0F4A3",x"10000",x"0F4C3",
									 x"10001",x"0FCE3",x"0FCE4",x"10001",x"0FD04",x"10008",x"0FD24",x"10010",x"0F504",x"10003",
									 x"0FD04",x"10003",x"0FCE4",x"0FCE3",x"10001",x"0FCC3",x"0F4A3",x"10001",x"0F483",x"0F463",
									 x"10000",x"0F462",x"0F442",x"10000",x"0F441",x"0F422",x"0F423",x"0EC23",x"0F444",x"0F466",
									 x"0F489",x"0F4EB",x"0F56F",x"0F5F3",x"0FE97",x"0FF1A",x"0FF9C",x"0FFDE",x"0FFFF",x"1004E",
									 x"0FFFF",x"1004C",x"0FFFE",x"0FF9C",x"0FF7B",x"0FF19",x"0FE95",x"0F632",x"0F58E",x"0ECCA",
									 x"0F467",x"0F426",x"0EC24",x"0EC43",x"0EC23",x"0EC22",x"0F442",x"0F462",x"10000",x"0F483",
									 x"10000",x"0F4A3",x"10000",x"0F4C3",x"0F4C4",x"10000",x"0FCE4",x"0FD04",x"0F4E4",x"0FD04",
									 x"10003",x"0FD24",x"10004",x"0FD44",x"10004",x"0FD64",x"10001",x"0FD44",x"10004",x"0FD64",
									 x"10000",x"0FD44",x"10008",x"0FD24",x"10004",x"0FD04",x"10002",x"0FCE4",x"10000",x"0F4E4",
									 x"0F4C4",x"10000",x"0F4A3",x"0F483",x"10000",x"0F462",x"10001",x"0F442",x"0F422",x"10000",
									 x"0F423",x"0F404",x"0F425",x"0EC67",x"0F4CA",x"0FD6D",x"0FDF1",x"0FE75",x"0FF19",x"0FF7C",
									 x"0FFBE",x"0FFDF",x"0FFFF",x"1004B",x"0FFFF",x"1004B",x"0FFBD",x"0FF5A",x"0FEB6",x"0FE33",
									 x"0F58F",x"0ECAA",x"0EC47",x"0EC25",x"0EC03",x"0EC23",x"0EC22",x"0EC42",x"10000",x"0F462",
									 x"10000",x"0F482",x"0F4A3",x"10000",x"0F4C3",x"10001",x"0F4E3",x"10000",x"0FCE4",x"0FD04",
									 x"10000",x"0FD25",x"0FD24",x"10000",x"0FD44",x"10004",x"0FD64",x"0FD65",x"0FD64",x"0FD44",
									 x"0FD64",x"0FD65",x"0FD64",x"10012",x"0FD65",x"0FD64",x"10002",x"0FD44",x"10004",x"0FD24",
									 x"10001",x"0FD04",x"10000",x"0FCE4",x"0F504",x"10001",x"0F4E4",x"10000",x"0F4C3",x"0FCC3",
									 x"0FCA3",x"10000",x"0FC83",x"0FC62",x"0FC42",x"0F442",x"0F402",x"10001",x"0F403",x"0F425",
									 x"0EC66",x"0ECA9",x"0F54E",x"0F613",x"0FEB7",x"0FF5A",x"0FFBD",x"0FFDF",x"0FFFF",x"10049",
									 x"0FFFF",x"10049",x"0FFBD",x"0FF5B",x"0F6F9",x"0F634",x"0F58F",x"0F50B",x"0EC88",x"0EC25",
									 x"0F403",x"10000",x"0EC02",x"0F422",x"0F442",x"0F462",x"10000",x"0F483",x"0F4A3",x"10000",
									 x"0F4C3",x"10000",x"0FCE3",x"0FCE4",x"10000",x"0FD04",x"10001",x"0FD24",x"10000",x"0FD45",
									 x"0FD24",x"0FD44",x"0FD45",x"10000",x"0FD44",x"10000",x"0FD64",x"10000",x"0FD65",x"0FD85",
									 x"0FD65",x"10001",x"0FD85",x"0FD65",x"0FD64",x"10008",x"0FD84",x"10001",x"0FD64",x"0F564",
									 x"0FD64",x"10000",x"0FD65",x"0FD64",x"0FD84",x"0FD85",x"0FD65",x"10001",x"0FD85",x"0FD65",
									 x"0FD64",x"10002",x"0FD45",x"10001",x"0FD25",x"0FD24",x"10002",x"0FD04",x"10001",x"0FCE3",
									 x"0F4E3",x"10000",x"0F4C3",x"10000",x"0F4A3",x"0F483",x"10000",x"0F463",x"0F462",x"0F442",
									 x"0F422",x"10000",x"0F424",x"0EC25",x"0F487",x"0F50A",x"0F58E",x"0F632",x"0FED7",x"0FF3B",
									 x"0FF9D",x"0FFDF",x"0FFFF",x"10047",x"0FFFF",x"10046",x"0FFDE",x"10000",x"0FF7C",x"0FED8",
									 x"0FE54",x"0F5D1",x"0ECEC",x"0EC47",x"0EC25",x"0EC24",x"0EC23",x"0F423",x"0F443",x"10000",
									 x"0F463",x"0FC83",x"0F4A3",x"10000",x"0FCA3",x"0FCC3",x"0F4C3",x"0F4E3",x"10000",x"0FD04",
									 x"10001",x"0FD24",x"10001",x"0FD45",x"10002",x"0FD65",x"10001",x"0FD64",x"10000",x"0FD84",
									 x"0FD85",x"10000",x"0FD84",x"0FD64",x"10001",x"0FD85",x"10000",x"0FDA5",x"0FD85",x"10001",
									 x"0FD86",x"10003",x"0FDA6",x"10001",x"0F5A6",x"10001",x"0FD86",x"0FD85",x"10003",x"0FD84",
									 x"0FD64",x"10001",x"0FD85",x"10000",x"0FD84",x"0FD64",x"10005",x"0FD44",x"10001",x"0FD24",
									 x"10001",x"0FD04",x"0F503",x"0F4E3",x"10001",x"0FCE4",x"0F4C3",x"0F4A4",x"10000",x"0F483",
									 x"10000",x"0F463",x"0F443",x"0F423",x"0F403",x"0F424",x"0EC25",x"0E467",x"0E4CA",x"0F5AF",
									 x"0FE34",x"0FEB8",x"0FF7C",x"0FFDD",x"0FFFF",x"10046",x"0FFFF",x"10045",x"0FFBE",x"0FF5B",
									 x"0FEF8",x"0FE54",x"0F56E",x"0F4CA",x"0F467",x"0F425",x"0F403",x"0F402",x"0F422",x"0F443",
									 x"0F463",x"0F483",x"10000",x"0FCA3",x"10000",x"0FCC4",x"10000",x"0FCE4",x"10000",x"0FD04",
									 x"0FD24",x"10001",x"0FD44",x"10002",x"0FD65",x"10002",x"0FD85",x"10001",x"0FD84",x"10001",
									 x"0FD85",x"0F585",x"10000",x"0FD64",x"0FD85",x"10000",x"0FDA6",x"0FDC7",x"0FDE8",x"0FE09",
									 x"10000",x"0FE2A",x"0FE0A",x"0FE2B",x"10000",x"0FE2C",x"10004",x"0FE2B",x"10001",x"0FE2A",
									 x"10000",x"0FE09",x"0FDE9",x"0FDE8",x"0FDC7",x"0FDA6",x"0FD85",x"0FD64",x"0FD85",x"10002",
									 x"0FD84",x"10000",x"0FD85",x"10000",x"0FD65",x"10002",x"0FD64",x"10000",x"0FD44",x"10002",
									 x"0FD24",x"0FD23",x"0FD24",x"10000",x"0FD04",x"0F4E4",x"10000",x"0F4C4",x"0F4C3",x"0F4A3",
									 x"10000",x"0F463",x"0F443",x"0F423",x"0F422",x"0F402",x"0EC03",x"0F424",x"0F467",x"0F4A9",
									 x"0F52E",x"0F633",x"0FEF8",x"0FF7B",x"0FFBE",x"0FFFF",x"10044",x"0FFFF",x"1003F",x"0F7DF",
									 x"0F7FF",x"0FFFF",x"10000",x"0FFDE",x"0FFBD",x"0FEF8",x"0FE74",x"0FDF1",x"0F50B",x"0EC46",
									 x"0EBE3",x"0F3E3",x"0F403",x"0F422",x"0F442",x"0F463",x"0F483",x"0F4A3",x"10000",x"0FCC4",
									 x"0FCE4",x"10001",x"0FD04",x"10001",x"0FD24",x"0FD44",x"10000",x"0FD45",x"0FD64",x"10001",
									 x"0FD65",x"10000",x"0FD64",x"0FD63",x"0FD83",x"0FD84",x"0FDA4",x"0FDA5",x"0FDA6",x"10000",
									 x"0FDC7",x"0FDE8",x"10001",x"0FE0A",x"0FE2A",x"0FE2B",x"0FE4D",x"0FE6E",x"0FE8F",x"0FE90",
									 x"10000",x"0FEB1",x"10000",x"0FED2",x"10000",x"0FED3",x"10004",x"0FED2",x"10001",x"0FEB1",
									 x"10000",x"0FEB0",x"0FE8F",x"0FE6F",x"0FE6E",x"0FE4C",x"0FE2B",x"0F60A",x"0FE09",x"0FDE8",
									 x"10000",x"0FDE7",x"10000",x"0FDC6",x"0FDA6",x"10000",x"0FD85",x"0FD65",x"10001",x"0FD64",
									 x"0FD84",x"0FD64",x"10002",x"0FD44",x"10000",x"0FD24",x"10001",x"0FD04",x"0F504",x"10000",
									 x"0F4E4",x"0F4C4",x"0F4C3",x"0F4A3",x"0F483",x"10000",x"0F442",x"0F422",x"0FC22",x"0FC03",
									 x"0F402",x"0F3E3",x"0EC26",x"0ECEB",x"0F5D0",x"0FE75",x"0FEF9",x"0F77C",x"0FFDE",x"0FFFF",
									 x"10042",x"0FFFF",x"10042",x"0FFDD",x"0FF5B",x"0FED6",x"0F5D0",x"0F50C",x"0F4A9",x"0EC46",
									 x"0F423",x"0F422",x"0F423",x"0F443",x"0F463",x"0F483",x"0F4A3",x"10000",x"0F4C3",x"0F4E4",
									 x"0FCE4",x"0FD04",x"10001",x"0FD24",x"0FD44",x"10000",x"0FD64",x"10000",x"0FD65",x"10000",
									 x"0FD64",x"0FD84",x"10000",x"0FD85",x"0FD65",x"10000",x"0FD84",x"10000",x"0F5A5",x"0F5C6",
									 x"0FDC8",x"0FDEA",x"0FE0B",x"0FE2C",x"0FE6E",x"10000",x"0FE8F",x"0FED1",x"0FEF2",x"0FF14",
									 x"0FF15",x"0FF36",x"10000",x"0FF37",x"10002",x"0FF58",x"10008",x"0FF38",x"0FF37",x"10002",
									 x"0FF36",x"10000",x"0FF15",x"0FF14",x"0FEF3",x"0FED1",x"0FEAF",x"0FE8E",x"0FE8D",x"0FE6C",
									 x"0F62B",x"0F608",x"0F5E7",x"0F5C6",x"0FDA5",x"0FD84",x"0FDA3",x"0FD84",x"0F565",x"0FD65",
									 x"10000",x"0FD84",x"10000",x"0FD64",x"10001",x"0FD44",x"10000",x"0FD24",x"10001",x"0F524",
									 x"0F504",x"0F4E4",x"0F4E3",x"0F4E4",x"0F4C4",x"0F4A3",x"0F463",x"10000",x"0F443",x"0F422",
									 x"10000",x"0F403",x"0EC45",x"0F4A8",x"0F50C",x"0F5B0",x"0FE96",x"0FF5A",x"0FFBD",x"0FFFF",
									 x"10041",x"0FFFF",x"1003F",x"0FFDE",x"0FFDD",x"0FF7B",x"0FE96",x"0F612",x"0FD6D",x"0F4A8",
									 x"0F425",x"0EC04",x"0EC23",x"0F441",x"0F462",x"0F463",x"0F483",x"0F4A4",x"0F4A3",x"0FCC3",
									 x"10000",x"0F4E3",x"0FD04",x"10000",x"0FD24",x"10001",x"0FD44",x"10000",x"0FD64",x"0FD85",
									 x"10000",x"0FD65",x"10000",x"0FD84",x"0F583",x"0FD84",x"0FDA5",x"0FDA7",x"0FDC9",x"0FDE9",
									 x"0FE0A",x"0FE2B",x"0FE4D",x"0FE8F",x"0FE91",x"0FEB2",x"0FEF4",x"0FEF5",x"0FF16",x"0FF36",
									 x"0FF57",x"0FF58",x"0FF79",x"0FF7A",x"10000",x"0FF7B",x"0FF7A",x"10000",x"0FF9A",x"10001",
									 x"0FFBA",x"0FF9A",x"0FF7A",x"0FF9A",x"10008",x"0FF7A",x"10003",x"0FF79",x"0FF58",x"0FF37",
									 x"0FF16",x"0FF15",x"0FEF4",x"0FED3",x"0FEB1",x"0FE8F",x"0FE4D",x"0FE2C",x"0FE0A",x"0FDE9",
									 x"0FDC8",x"0FDA7",x"0FDA6",x"0FD85",x"0FD84",x"10000",x"0FD85",x"10001",x"0FD64",x"10000",
									 x"0FD44",x"10000",x"0F544",x"0F524",x"10000",x"0F504",x"0FD04",x"0FCE3",x"10000",x"0FCC3",
									 x"0F4A3",x"10001",x"0F483",x"0EC63",x"0F443",x"0F402",x"10000",x"0F425",x"0F488",x"0F54D",
									 x"0FE12",x"0FE96",x"0FF5B",x"0FFBD",x"0FFDE",x"0FFFF",x"1003E",x"0FFFF",x"1003C",x"0FFDE",
									 x"10000",x"0FFBD",x"0FF5B",x"0FEF8",x"0F613",x"0ED0C",x"0F4A8",x"0F445",x"0EC03",x"0F423",
									 x"0F422",x"0F462",x"0F482",x"0FCA3",x"0F483",x"0F4A3",x"0FCE4",x"10000",x"0FCE3",x"0FD03",
									 x"0FD24",x"10000",x"0FD45",x"0FD65",x"0FD64",x"10000",x"0FD85",x"10000",x"0FD65",x"0FD85",
									 x"10001",x"0FDA5",x"0FDC6",x"0FDE7",x"0F609",x"0F62B",x"0FE4E",x"0FE71",x"0FEB2",x"0FEF3",
									 x"0FF15",x"0FF36",x"0FF58",x"0FF79",x"10001",x"0FF9A",x"10000",x"0FF7A",x"0FF79",x"10000",
									 x"0FF7A",x"0FF9A",x"1001B",x"0FF99",x"10002",x"0FF79",x"0FF78",x"0FF57",x"0FF15",x"0FEF3",
									 x"0FED2",x"0FE8F",x"0FE6E",x"0F62C",x"0F5E9",x"0FDC8",x"0FDC6",x"0FDA6",x"0FD85",x"0FD84",
									 x"10000",x"0FD85",x"0FD65",x"0FD64",x"10000",x"0FD44",x"10001",x"0FD24",x"10000",x"0FD04",
									 x"0FCE4",x"0FCE3",x"10000",x"0F4E3",x"0F4C3",x"0F483",x"10000",x"0F463",x"0F422",x"10000",
									 x"0EC03",x"0F445",x"0F488",x"0F50C",x"0FE12",x"0FEB7",x"0FF3B",x"0FFBD",x"0FFFF",x"1003D",
									 x"0FFFF",x"1003C",x"0FFDE",x"0FFBD",x"0FEF9",x"0EE34",x"0ED6F",x"0ECAA",x"0EC26",x"0F404",
									 x"0F403",x"0F423",x"0F463",x"0F483",x"0F4A3",x"0FCC3",x"10001",x"0FCE4",x"0FD04",x"0FD24",
									 x"10000",x"0FD44",x"0FD45",x"0FD65",x"10000",x"0FD85",x"10004",x"0FDA5",x"0F5A5",x"0F5C6",
									 x"0FE08",x"0FE4B",x"0FE8E",x"0FEB1",x"0FEF3",x"0FF35",x"0FF57",x"0FF78",x"10000",x"0FF79",
									 x"0FF9A",x"10006",x"0FF7A",x"10001",x"0FF79",x"10001",x"0FF7A",x"0FF9A",x"1001B",x"0FF9B",
									 x"10000",x"0FF9A",x"0FF79",x"0FF78",x"0FF77",x"0FF76",x"0FF55",x"0FF13",x"0FED0",x"0FE8E",
									 x"0FE2C",x"0FDE9",x"0FDA7",x"0FDA6",x"0FDA5",x"0FD85",x"0FD64",x"0FD84",x"10000",x"0FD85",
									 x"0FD65",x"10000",x"0FD44",x"10000",x"0FD24",x"10000",x"0FD04",x"0FD03",x"0F503",x"0F4E3",
									 x"0FCC3",x"0F4A3",x"0F483",x"0F463",x"0F442",x"0F422",x"0F423",x"0F403",x"0E405",x"0E4AA",
									 x"0ED4F",x"0F613",x"0F6F8",x"0FF9D",x"0FFDE",x"0FFFF",x"1003B",x"0FFFF",x"10038",x"0FFFE",
									 x"0FFFF",x"10000",x"0FFDF",x"0FF9C",x"0FF3A",x"0FE33",x"0F54D",x"0F4A9",x"0F425",x"0F3E3",
									 x"0F403",x"0F423",x"0F443",x"0F463",x"0F483",x"0F4A3",x"0F4C3",x"0FCE4",x"0FD04",x"10000",
									 x"0FD24",x"10000",x"0FD44",x"0F544",x"0F565",x"0FD65",x"10000",x"0FD85",x"0FD84",x"10000",
									 x"0FD85",x"10000",x"0F5A6",x"0F5E7",x"0F628",x"0F62B",x"0FE6E",x"0FEB1",x"0FEF4",x"0FF17",
									 x"0FF39",x"0FF7A",x"0FF9A",x"10006",x"0FF7A",x"10003",x"0FF79",x"10000",x"0FF99",x"10010",
									 x"0FF9A",x"0FF99",x"10006",x"0FF79",x"10004",x"0FF7A",x"0FF9B",x"0FF9A",x"0FF7A",x"10000",
									 x"0FF9A",x"0FF7A",x"0FF79",x"0FF58",x"0FF36",x"0FEF4",x"0FEB2",x"0FE6F",x"0FE2C",x"0F5EA",
									 x"0FDE8",x"0FDA6",x"0FD85",x"0FD84",x"0F584",x"0FD85",x"10000",x"0FD65",x"0FD85",x"0FD65",
									 x"0FD44",x"10000",x"0FD24",x"10000",x"0F504",x"10000",x"0FCE3",x"0F4C3",x"0F4A3",x"0F483",
									 x"10000",x"0F462",x"0F422",x"0F402",x"0EBE2",x"0EC25",x"0F4A8",x"0F52C",x"0FE12",x"0FF18",
									 x"0FF9D",x"0FFDE",x"0FFFF",x"1003A",x"0FFFF",x"10039",x"0FFDF",x"0FFBE",x"0FF3A",x"0FE95",
									 x"0F5AF",x"0ECCA",x"0EC26",x"0F403",x"0FC02",x"0F422",x"0F463",x"10000",x"0F483",x"0F4A3",
									 x"0F4C3",x"0FCE3",x"0FD04",x"0F504",x"0FD24",x"0FD44",x"10000",x"0FD64",x"10001",x"0FD65",
									 x"10001",x"0FD85",x"0FDA5",x"0FDC6",x"0FDC7",x"0FDE9",x"0FE4C",x"0FE8F",x"0FED1",x"0FEF4",
									 x"0FF16",x"0FF37",x"0FF58",x"0FF59",x"0FF7A",x"10002",x"0FF9A",x"0FF7A",x"10001",x"0FF9A",
									 x"10001",x"0FF7A",x"10002",x"0FF9A",x"0FF99",x"10002",x"0FF9A",x"0FF99",x"10013",x"0FF79",
									 x"10006",x"0FF99",x"0FF9A",x"10003",x"0FF9B",x"0FF7A",x"10000",x"0FF79",x"0FF78",x"0FF58",
									 x"0FF56",x"0FF15",x"0FED2",x"0FE8F",x"0FE4C",x"0FE0A",x"0FDE8",x"0FDA6",x"0FDA5",x"0FD85",
									 x"10001",x"0FD84",x"0FD64",x"0FD44",x"10000",x"0FD24",x"0FD25",x"0F524",x"0FD04",x"10000",
									 x"0FCE4",x"0FCC4",x"0F4A3",x"0F483",x"0F463",x"0F442",x"10000",x"0EC23",x"0EC43",x"0EC24",
									 x"0EC88",x"0ED8F",x"0F676",x"0FF1A",x"0FF9D",x"0FFDF",x"10000",x"0FFFF",x"10037",x"0FFFF",
									 x"10038",x"0F7DE",x"0FF7C",x"0FEB7",x"0F5B1",x"0F4EB",x"0EC66",x"0EC24",x"0EC03",x"0F423",
									 x"0FC42",x"0F483",x"0F4A3",x"0F4C4",x"0FCC4",x"0FCE4",x"0FD04",x"0FD24",x"10002",x"0FD44",
									 x"0FD65",x"0FD84",x"0FDA5",x"10001",x"0FD85",x"0FD86",x"0FDA7",x"0FDE9",x"0FE4C",x"0FE8E",
									 x"0FED1",x"0FF14",x"0FF37",x"0FF39",x"0FF5A",x"0FF7A",x"10000",x"0FF99",x"10002",x"0FF79",
									 x"10001",x"0FF99",x"10001",x"0FF9A",x"10001",x"0FF7A",x"10000",x"0FF79",x"10000",x"0FF99",
									 x"1001C",x"0FF79",x"10003",x"0FF99",x"10003",x"0FF9A",x"10002",x"0FF99",x"10001",x"0FF9A",
									 x"0FF79",x"0FF58",x"0FF56",x"0FF14",x"0FEF2",x"0FEAF",x"0FE4C",x"0FDE9",x"0FDA7",x"0FD86",
									 x"0FD85",x"0F585",x"0FD84",x"0FD85",x"0FD65",x"0FD45",x"0FD65",x"0F545",x"0FD24",x"0F524",
									 x"0FD04",x"10000",x"0FCE4",x"0F4C4",x"0F4C3",x"0F4A3",x"0F483",x"0F442",x"0EC22",x"10000",
									 x"0EC24",x"0E467",x"0E50C",x"0EDB0",x"0FE96",x"0FF5B",x"0FF9D",x"0FFDE",x"0FFFF",x"10036",
									 x"0FFFF",x"10037",x"0FFDE",x"0FF5B",x"0FEB6",x"0FDB0",x"0F4AA",x"0F446",x"0EC04",x"0F422",
									 x"10000",x"0FC63",x"0FC83",x"0F4C2",x"10000",x"0F4E3",x"0F4E4",x"0F504",x"10000",x"0FD44",
									 x"0FD45",x"10000",x"0FD44",x"0FD65",x"0FD64",x"0FD84",x"10000",x"0FDA5",x"0FDC6",x"0FDC7",
									 x"0FDC9",x"0F60B",x"0FE6E",x"0FEB2",x"0FF15",x"0FF57",x"0FF98",x"0FF79",x"0FF7A",x"10002",
									 x"0FF79",x"10003",x"0FF99",x"10001",x"0FF9A",x"10000",x"0FF99",x"10028",x"0FF7A",x"10000",
									 x"0FF79",x"10004",x"0FF99",x"0FF79",x"10000",x"0FF9A",x"10000",x"0FF7A",x"10001",x"0FF79",
									 x"0FF57",x"0FF35",x"0FED3",x"0FE6F",x"0FE0B",x"0FDC9",x"0F5C8",x"0F5A6",x"0FDA5",x"0FD85",
									 x"10000",x"0FD65",x"0FD85",x"0F565",x"0FD44",x"10000",x"0FD24",x"0F504",x"10000",x"0F4E3",
									 x"10001",x"0F4C3",x"0F4A3",x"0F462",x"0F442",x"0F402",x"0EC03",x"0EC45",x"0F4A9",x"0F5AF",
									 x"0FE96",x"0FF3A",x"0FFBC",x"0FFFE",x"0FFFF",x"10035",x"0FFFF",x"10036",x"0FFBE",x"0F739",
									 x"0F633",x"0F54E",x"0F4A9",x"0FC25",x"0F403",x"0EC43",x"0F442",x"0F462",x"0F483",x"0F4C3",
									 x"0F4E3",x"10000",x"0F503",x"0F523",x"0FD24",x"0F524",x"0FD44",x"0FD65",x"10002",x"0FD84",
									 x"0FD85",x"0FD86",x"0FDC7",x"0FDE9",x"0FE2C",x"0FE8F",x"0FED2",x"0FF14",x"0FF37",x"0FF79",
									 x"0FF99",x"10001",x"0FF79",x"10002",x"0FF59",x"0FF79",x"10003",x"0FF99",x"10002",x"0FF79",
									 x"10003",x"0FF99",x"0FF79",x"10004",x"0FF99",x"1001C",x"0FF79",x"1000D",x"0FF9A",x"10000",
									 x"0FF79",x"0FF58",x"0FF57",x"0FF15",x"0FED2",x"0FE90",x"0F62C",x"0F5E9",x"0F5C7",x"0FDA5",
									 x"0FD85",x"10001",x"0F565",x"0F564",x"0F565",x"0F545",x"0F544",x"0F524",x"0F523",x"0FD03",
									 x"0F4E3",x"0FCC3",x"10000",x"0F4A3",x"0F483",x"0F442",x"0EC22",x"0F422",x"0EC24",x"0F4A8",
									 x"0FD4D",x"0F613",x"0FF19",x"0FFBE",x"0FFFF",x"10035",x"0FFFF",x"10032",x"0FFDF",x"0FFFF",
									 x"0FFBE",x"0FF5C",x"0FED8",x"0EDF2",x"0E50B",x"0E468",x"0EC04",x"0F403",x"0F443",x"0F483",
									 x"10000",x"0F4A4",x"0FCC4",x"0F4E3",x"0FD04",x"0FD03",x"0F523",x"0FD24",x"0FD45",x"0FD65",
									 x"10000",x"0FD85",x"10002",x"0FDA5",x"0FDC7",x"0FE09",x"0FE4C",x"0FE8F",x"0FEF2",x"0FF55",
									 x"0FF77",x"0FF98",x"0FF99",x"10000",x"0FF79",x"10007",x"0FF99",x"10000",x"0FF79",x"10013",
									 x"0FF99",x"1001A",x"0FF79",x"1000B",x"0FF99",x"10000",x"0FF79",x"10001",x"0FF99",x"0FF79",
									 x"0FF78",x"0FF56",x"0FEF3",x"0FEB0",x"0FE6C",x"0FE0A",x"0FDE7",x"0FDC6",x"0FDA5",x"0FD85",
									 x"0FD84",x"0FD85",x"0FD65",x"10000",x"0FD64",x"0FD44",x"0FD24",x"0FD04",x"10000",x"0FCE4",
									 x"0F4C3",x"10000",x"0F483",x"0F462",x"0F442",x"0EC23",x"0EC04",x"0EC46",x"0E4CA",x"0EDD1",
									 x"0F6D9",x"0F75B",x"0FFBD",x"0FFFE",x"0FFFF",x"10032",x"0FFFF",x"10033",x"0FFDE",x"0FF3A",
									 x"0FE96",x"0FDB1",x"0ECCA",x"0EC45",x"0EC23",x"0F442",x"0F462",x"0FC82",x"0FCA3",x"0F4A3",
									 x"0F4C4",x"0FCE4",x"0FD04",x"0FD24",x"10000",x"0FD44",x"0FD45",x"0FD65",x"10001",x"0FD85",
									 x"0FD84",x"0FDA4",x"0FDC6",x"0FE09",x"0FE4C",x"0FEAF",x"0FEF3",x"0FF36",x"0FF98",x"0FF99",
									 x"10000",x"0FF7A",x"0FF79",x"10009",x"0FF99",x"10000",x"0FF79",x"1002B",x"0FF99",x"10002",
									 x"0FF79",x"10010",x"0FF9A",x"10000",x"0FF7A",x"0FF79",x"0FF77",x"0FF56",x"0FF14",x"0FEB0",
									 x"0FE4C",x"0FE09",x"0FDC7",x"0FDA5",x"0FDA4",x"0FD84",x"10000",x"0FD65",x"0FD64",x"0FD44",
									 x"10000",x"0FD24",x"10000",x"0FD04",x"0FCE4",x"10000",x"0F4C3",x"0F483",x"0F462",x"0F442",
									 x"0F423",x"0EC03",x"0E404",x"0E489",x"0F58F",x"0FE54",x"0FF39",x"0FFDE",x"0FFFF",x"10032",
									 x"0FFFF",x"10031",x"0FFDE",x"0FFBE",x"0FF5A",x"0FE54",x"0FD6E",x"0FCA9",x"0F424",x"0F3E2",
									 x"0F422",x"0F442",x"0F482",x"0F4A3",x"0FCC3",x"0FCE4",x"0FD04",x"10000",x"0FD24",x"0FD44",
									 x"0FD64",x"0FD65",x"10000",x"0FD64",x"10000",x"0FD84",x"0FD85",x"0FDC6",x"0FDE7",x"0FE2B",
									 x"0FE6F",x"0FED3",x"0FF15",x"0FF58",x"0FF79",x"0FF99",x"10000",x"0FF79",x"10007",x"0FF78",
									 x"10000",x"0FF79",x"10000",x"0FF99",x"10000",x"0FF79",x"10009",x"0FF99",x"0FF79",x"1001F",
									 x"0FF99",x"10002",x"0FF79",x"10006",x"0FF99",x"10000",x"0FF79",x"10008",x"0FF7A",x"0FF79",
									 x"10001",x"0FF59",x"0FF16",x"0FED2",x"0FE6E",x"0FE2B",x"0FDE8",x"0FDC6",x"0FDA5",x"0FD85",
									 x"0FD65",x"10001",x"0FD64",x"0FD44",x"10000",x"0FD24",x"0FD04",x"10000",x"0F4E4",x"0F4C3",
									 x"0F4A3",x"0F483",x"0F463",x"0F422",x"0F402",x"0F424",x"0FCA9",x"0FD2D",x"0FE34",x"0FF3B",
									 x"0FFBE",x"0FFDF",x"0FFFF",x"10030",x"0FFFF",x"10030",x"0FFDE",x"0FF7C",x"0FEF9",x"0F633",
									 x"0ED0B",x"0EC26",x"0EBE3",x"0F402",x"0FC22",x"0FC43",x"0F483",x"0F4C3",x"0FCE4",x"10000",
									 x"0FD04",x"0FD24",x"10000",x"0FD44",x"0FD65",x"0FD85",x"10000",x"0FD84",x"0FDA4",x"10000",
									 x"0FDC6",x"0FDE7",x"0FE2B",x"0FE6E",x"0FEB1",x"0FF15",x"0FF38",x"0FF5A",x"0FF7A",x"0FF79",
									 x"10000",x"0FF78",x"1000C",x"0FF98",x"10000",x"0FF78",x"1000A",x"0FF79",x"1000A",x"0FF78",
									 x"1001F",x"0FF98",x"10000",x"0FF78",x"10002",x"0FF79",x"10000",x"0FF78",x"10000",x"0FF58",
									 x"10001",x"0FF79",x"10001",x"0FF7A",x"0FF79",x"0FF57",x"0FF34",x"0FEB0",x"0FE6E",x"0FE2B",
									 x"0FDE8",x"0FDC6",x"0FD85",x"10001",x"0FD84",x"0FD64",x"10000",x"0FD44",x"0FD24",x"10000",
									 x"0F504",x"0F4E3",x"10000",x"0F4C3",x"0F483",x"0F442",x"0FC22",x"0F403",x"0EBE4",x"0F427",
									 x"0ECEC",x"0FE14",x"0FEF9",x"0FF7C",x"0FFDE",x"0FFFF",x"1002F",x"0FFFF",x"1002F",x"0FFDE",
									 x"0FF7C",x"0F6B7",x"0F5F2",x"0ED0C",x"0EC46",x"0F3E3",x"0F402",x"0F462",x"0FC83",x"10000",
									 x"0FCC4",x"10000",x"0F504",x"0FD04",x"0FD24",x"0FD44",x"0FD64",x"10000",x"0FD85",x"10001",
									 x"0FDA5",x"10000",x"0FDC6",x"0FE09",x"0FE4C",x"0FEB0",x"0FEF3",x"0FF36",x"0FF58",x"0FF79",
									 x"0FF59",x"0FF79",x"10000",x"0FF78",x"10001",x"0FF58",x"10000",x"0FF78",x"10016",x"0FF79",
									 x"1000A",x"0FF78",x"1001F",x"0FF98",x"0FF78",x"10003",x"0FF79",x"10000",x"0FF78",x"0FF79",
									 x"0FF59",x"10000",x"0FF58",x"10000",x"0FF78",x"10000",x"0FF79",x"10001",x"0FF78",x"0FF36",
									 x"0FEF4",x"0FEB1",x"0FE4D",x"0FE09",x"0FDC6",x"0FDA5",x"10000",x"0FD84",x"10001",x"0FD64",
									 x"0FD44",x"10000",x"0FD24",x"0F504",x"10000",x"0F4E4",x"0F4C3",x"0F4A3",x"0FCA2",x"0F463",
									 x"0F403",x"10000",x"0EC25",x"0F4EB",x"0F5D1",x"0FE97",x"0FF5C",x"0FFDF",x"0FFFF",x"1002E",
									 x"0FFFF",x"1002E",x"0FFDF",x"0FFBD",x"0FEF8",x"0F5D1",x"0F4EB",x"0EC67",x"0EC04",x"0F423",
									 x"0F443",x"0F483",x"0F4A3",x"10000",x"0FCC3",x"0FCE4",x"0FD04",x"0FD24",x"0FD44",x"0FD64",
									 x"10000",x"0FD84",x"0F584",x"0F5A3",x"0F584",x"0FD85",x"0FDC7",x"0FDE9",x"0FE4D",x"0FEB1",
									 x"0FF15",x"0FF57",x"0FF78",x"10009",x"0FF58",x"10000",x"0FF78",x"1004B",x"0FF79",x"0FF78",
									 x"0FF58",x"10003",x"0FF78",x"0FF58",x"10001",x"0FF57",x"0FF35",x"0FED2",x"0FE4D",x"0FE09",
									 x"0FDC7",x"0FDA5",x"0FDA4",x"0F5A3",x"0F5A4",x"0FDA4",x"0FD85",x"0FD64",x"0FD44",x"0F524",
									 x"0F504",x"10000",x"0F4E4",x"0F4C3",x"10000",x"0F483",x"0F442",x"0F423",x"0EC02",x"0F465",
									 x"0ECCA",x"0F5B1",x"0F6B8",x"0FF9D",x"0FFDE",x"0FFFF",x"1002D",x"0FFFF",x"1002D",x"0FFDE",
									 x"0FF7B",x"0FEF8",x"0EDD1",x"0ECA9",x"0EC25",x"0EC04",x"0F443",x"0F462",x"0F483",x"0F4C3",
									 x"0FCE4",x"10000",x"0FD04",x"10001",x"0FD25",x"0FD45",x"0FD65",x"0FD85",x"10000",x"0F5A4",
									 x"0FDA4",x"0FDA5",x"0FDC8",x"0FE0C",x"0FE8F",x"0FEF2",x"0FF36",x"0FF58",x"10000",x"0FF78",
									 x"10003",x"0FF58",x"10000",x"0FF78",x"10000",x"0FF58",x"0FF78",x"10051",x"0FF58",x"10005",
									 x"0FF78",x"10001",x"0FF56",x"0FED3",x"0FE8F",x"0FE4B",x"0FDE9",x"0FDA6",x"0FDA4",x"0FDC4",
									 x"0FDA5",x"10000",x"0FD84",x"0FD64",x"0FD44",x"10000",x"0FD24",x"0FD04",x"0F4E4",x"0F4C4",
									 x"0F4A3",x"0F483",x"0F463",x"0EC22",x"0F422",x"0EC04",x"0E489",x"0ED90",x"0FEB7",x"0FF5B",
									 x"0FFDE",x"10000",x"0FFFF",x"1002B",x"0FFFF",x"1002C",x"0FFBE",x"0FF1A",x"0F613",x"0F58F",
									 x"0ECA9",x"0EC04",x"0F402",x"0F422",x"0FC62",x"0F482",x"0F4C2",x"0F4E3",x"0FD04",x"10000",
									 x"0FD24",x"0FD25",x"10000",x"0FD45",x"0FD46",x"0FD65",x"10000",x"0FD85",x"0FDA6",x"0FDC8",
									 x"0FE0A",x"0FE6F",x"0FED3",x"0FF15",x"0FF57",x"0FF58",x"10002",x"0FF78",x"10006",x"0FF58",
									 x"0FF78",x"10052",x"0FF58",x"10004",x"0FF78",x"0FF58",x"0FF59",x"0FF79",x"0FF58",x"0FF15",
									 x"0FEF3",x"0FE90",x"0FE0B",x"0FDC7",x"0FDA5",x"0FD85",x"0FD65",x"10000",x"0FD64",x"10000",
									 x"0FD65",x"0FD45",x"0FD24",x"0FD04",x"10000",x"0F4E4",x"0F4A3",x"10000",x"0F463",x"0F442",
									 x"0F3E2",x"0EC04",x"0EC68",x"0FD6E",x"0F613",x"0FF19",x"0FFBC",x"0FFFE",x"0FFFF",x"10000",
									 x"0FFDF",x"0FFFF",x"10027",x"0FFFF",x"10028",x"0FFFE",x"0FFFF",x"10000",x"0FFDF",x"0FF7D",
									 x"0FE76",x"0ED2D",x"0F4A8",x"0EC24",x"0F402",x"0FC42",x"0FC63",x"0FCA3",x"0FCC3",x"0FCE3",
									 x"0FD04",x"0FD24",x"10000",x"0FD44",x"0FD45",x"0FD65",x"10000",x"0FD85",x"0FD84",x"0FDA4",
									 x"0FDC5",x"0FDE7",x"0FE0A",x"0FE8E",x"0FEF3",x"0FF57",x"0FF79",x"10000",x"0FF59",x"0FF58",
									 x"0FF78",x"10002",x"0FF77",x"0FF78",x"10058",x"0FF77",x"0FF57",x"10002",x"0FF78",x"0FF57",
									 x"0FF58",x"10000",x"0FF59",x"0FF79",x"0FF78",x"0FF57",x"0FF15",x"0FE8F",x"0FE0A",x"0FDC7",
									 x"0FDA6",x"0FD85",x"10001",x"0FD64",x"0FD65",x"10000",x"0FD45",x"0FD24",x"10000",x"0F504",
									 x"0F4C4",x"10000",x"0FCA4",x"0F463",x"0FC42",x"0F423",x"0F404",x"0F467",x"0ED0C",x"0F634",
									 x"0FF7B",x"0FFDE",x"0FFFF",x"10000",x"0FFFE",x"0FFFF",x"10027",x"0FFFF",x"10029",x"0FFFE",
									 x"0FFDE",x"0FF7C",x"0FEB7",x"0F590",x"0EC88",x"0EC45",x"0EC23",x"0F422",x"0F442",x"0F463",
									 x"0F4C3",x"0F4E4",x"10000",x"0FD05",x"0FD24",x"0FD44",x"0FD45",x"0FD65",x"10000",x"0FD85",
									 x"0FDA4",x"10000",x"0FDC5",x"0F5E7",x"0FE4B",x"0FE8E",x"0FF12",x"0FF56",x"0FF78",x"10000",
									 x"0FF58",x"0FF38",x"0FF58",x"10000",x"0FF57",x"10000",x"0FF77",x"10060",x"0FF57",x"10001",
									 x"0FF78",x"10002",x"0FF57",x"0FF13",x"0FEAF",x"0FE4B",x"0FDE9",x"0FDA6",x"0FDA5",x"0F584",
									 x"0FD84",x"10000",x"0FD65",x"10000",x"0FD44",x"10000",x"0F524",x"0F4E3",x"10000",x"0FCC3",
									 x"0F483",x"0F463",x"0F443",x"0F402",x"0F404",x"0EC67",x"0ED4E",x"0FE96",x"0FF5C",x"0FFDF",
									 x"0FFFF",x"0FFFE",x"10000",x"0FFFF",x"10026",x"0FFFF",x"10029",x"0FFBD",x"0FF5A",x"0FEB6",
									 x"0F56E",x"0E447",x"0EBE4",x"0EC03",x"0F463",x"0FCA3",x"0FCC3",x"0F4C3",x"0F4E4",x"0F504",
									 x"0FD24",x"10000",x"0FD65",x"10000",x"0FD85",x"10002",x"0F5C5",x"0F5E6",x"0FDEA",x"0FE2E",
									 x"0FED2",x"0FF15",x"0FF56",x"0FF78",x"0FF58",x"0FF57",x"0FF56",x"0FF37",x"0FF58",x"0FF78",
									 x"0FF57",x"10000",x"0FF77",x"10060",x"0FF57",x"10000",x"0FF37",x"0FF57",x"0FF77",x"10000",
									 x"0FF78",x"10000",x"0FF57",x"0FF54",x"0FEF1",x"0FE6E",x"0F60A",x"0FDE6",x"0FDA5",x"0F584",
									 x"0FD85",x"10001",x"0FD65",x"0FD64",x"0FD44",x"0FD24",x"0FD04",x"0FCE4",x"0F4C3",x"0F4A4",
									 x"10000",x"0F463",x"0F402",x"0EC03",x"0EC66",x"0F54D",x"0FE75",x"0FF5B",x"0FFBD",x"0FFFE",
									 x"0FFFF",x"10027",x"0FFFF",x"10029",x"0FF5C",x"0F696",x"0ED8F",x"0EC88",x"0EC24",x"0F423",
									 x"0F422",x"0F483",x"0F4C3",x"10000",x"0F4E3",x"0F524",x"10000",x"0FD44",x"10000",x"0FD65",
									 x"0FD85",x"10003",x"0FDC7",x"0FE2A",x"0FE6F",x"0FEB3",x"0FF17",x"0FF38",x"0FF58",x"0FF57",
									 x"0FF37",x"10000",x"0FF36",x"0FF37",x"10000",x"0FF57",x"10002",x"0FF77",x"0FF57",x"0FF77",
									 x"1005D",x"0FF57",x"10000",x"0FF37",x"0FF36",x"0FF57",x"10000",x"0FF37",x"0FF57",x"0FF58",
									 x"0FF77",x"0FF56",x"0FEF3",x"0FE8F",x"0FE2A",x"0FDE6",x"0F5A5",x"10000",x"0FDA6",x"10000",
									 x"0FD85",x"10000",x"0FD64",x"0FD44",x"0FD24",x"0FD04",x"0FCE4",x"0F4C4",x"0F4A3",x"0F483",
									 x"0F442",x"0F422",x"0EC23",x"0EC87",x"0ED4D",x"0F675",x"0FF5B",x"0FFDE",x"0FFFF",x"10027",
									 x"0FFFF",x"10027",x"0FFDF",x"0FF9D",x"0FED7",x"0F5B0",x"0F4CA",x"0EC45",x"0EC23",x"0F442",
									 x"0F462",x"0F4A3",x"0F4E3",x"10000",x"0F504",x"0FD24",x"0F524",x"0FD45",x"0FD65",x"0FD84",
									 x"0FD85",x"10001",x"0FD86",x"0FDA6",x"0FE0A",x"0FE8E",x"0FED2",x"0FF15",x"0FF57",x"10010",
									 x"0FF77",x"1004E",x"0FF57",x"10000",x"0FF77",x"10003",x"0FF57",x"10009",x"0FF56",x"0FF57",
									 x"10000",x"0FF58",x"10000",x"0FF15",x"0FED2",x"0FE8F",x"0FE2A",x"0F5E7",x"0F5C5",x"0F5A6",
									 x"0FDA6",x"0FDA5",x"0FD85",x"0F564",x"0F544",x"0FD44",x"0FD24",x"0FD04",x"0F4E4",x"0F4C3",
									 x"0F4A3",x"0F462",x"0F442",x"0F422",x"0EC25",x"0ECA9",x"0F5B0",x"0FE96",x"0FF9C",x"0FFDE",
									 x"10000",x"0FFFF",x"10025",x"0FFFF",x"10026",x"0FFFE",x"0FF7B",x"0FEB7",x"0FD8F",x"0ECA8",
									 x"0EC45",x"0EC23",x"0F443",x"0FC82",x"0F483",x"0F4C4",x"0F504",x"10000",x"0FD24",x"0FD45",
									 x"10000",x"0FD65",x"0FD85",x"0FDA4",x"0FD84",x"10000",x"0FDA5",x"0FDC7",x"0FE0A",x"0FE90",
									 x"0FEF3",x"0FF35",x"0FF56",x"0FF57",x"10020",x"0FF77",x"10032",x"0FF57",x"1001C",x"0FF56",
									 x"0FF57",x"10002",x"0FF56",x"0FF35",x"0FF14",x"0FEB0",x"0FE4B",x"0FDE8",x"0FDA6",x"0FDA5",
									 x"10002",x"0FD65",x"10000",x"0FD45",x"0FD24",x"0F524",x"0F4E4",x"0F4C4",x"0F4A3",x"0F483",
									 x"0F463",x"0F423",x"0F424",x"0EC88",x"0F56E",x"0FEB6",x"0FF7B",x"0FFBD",x"0FFFF",x"10025",
									 x"0FFFF",x"10026",x"0F79B",x"0F6B7",x"0F590",x"0EC68",x"0EC04",x"0EC22",x"0F443",x"0FC83",
									 x"0FCA2",x"0F4C3",x"0F504",x"0F524",x"0FD24",x"0FD44",x"0FD65",x"10000",x"0FD85",x"0FDA5",
									 x"0FDC5",x"0FDA4",x"10000",x"0FDE7",x"0FE4B",x"0FECF",x"0FF15",x"0FF37",x"0FF57",x"0FF37",
									 x"0FF57",x"0FF56",x"10000",x"0FF57",x"0FF56",x"0FF57",x"10001",x"0FF56",x"10008",x"0FF57",
									 x"10003",x"0FF56",x"10008",x"0FF57",x"10000",x"0FF77",x"10030",x"0FF57",x"10000",x"0FF56",
									 x"1000A",x"0FF57",x"10002",x"0FF56",x"0FF57",x"0FF56",x"10001",x"0FF57",x"10000",x"0FF56",
									 x"10005",x"0FF57",x"10000",x"0FF56",x"10001",x"0FF57",x"0FF58",x"0FF35",x"0FEB0",x"0FE2B",
									 x"0FDE8",x"0FDA6",x"0FDA5",x"10000",x"0FDC5",x"0FD85",x"10000",x"0FD65",x"0FD44",x"0FD24",
									 x"0F504",x"0FD04",x"0F4C4",x"0F4A3",x"0F483",x"0F443",x"0F402",x"0F403",x"0EC88",x"0ED8F",
									 x"0F696",x"0FF5A",x"0FFDE",x"0FFFF",x"10024",x"0FFFF",x"10024",x"0FFDF",x"0FFBD",x"0F718",
									 x"0F612",x"0F4EB",x"0EC25",x"0EC23",x"0EC42",x"0F463",x"0F4A2",x"0F4C3",x"0F4E4",x"0F504",
									 x"0F524",x"0FD44",x"0FD64",x"10000",x"0FD85",x"0F584",x"0FDA5",x"10000",x"0F5A5",x"0F5E7",
									 x"0FE2B",x"0FE8F",x"0FF13",x"0FF36",x"0FF57",x"10001",x"0FF56",x"10000",x"0FF36",x"0FF56",
									 x"10075",x"0FF57",x"0FF58",x"0FF57",x"0FF14",x"0FE90",x"0FE2C",x"0FDC8",x"0FDA5",x"10002",
									 x"0FD85",x"0FD65",x"0FD64",x"0FD44",x"0FD24",x"0F504",x"0F4E4",x"0F4E3",x"0F4A3",x"0F483",
									 x"0EC22",x"0F402",x"0EC25",x"0E4CA",x"0F5F1",x"0F6D6",x"0FF9C",x"0FFFF",x"0F7FF",x"0FFFF",
									 x"10022",x"0FFFF",x"10023",x"0FFDF",x"0FFBD",x"0FF3A",x"0FDF2",x"0F50C",x"0F466",x"0F422",
									 x"0F442",x"0EC63",x"0F4A4",x"0F4C3",x"0F4E3",x"0FD04",x"0FD25",x"0FD44",x"0FD64",x"10000",
									 x"0FD84",x"0FDA5",x"0FDA4",x"0FDA5",x"0FDC5",x"0FDE7",x"0F64C",x"0FEB0",x"0FF14",x"0FF36",
									 x"10001",x"0FF56",x"10077",x"0FF36",x"10001",x"0FF56",x"10001",x"0FF55",x"0FF14",x"0FEB1",
									 x"0FE2C",x"0FDE7",x"0FDC5",x"0FDA5",x"10001",x"0FD85",x"10000",x"0FD64",x"0FD44",x"0FD24",
									 x"0F504",x"0FD04",x"0F4E3",x"0F4A3",x"0F462",x"0F422",x"0F424",x"0EC46",x"0F4EA",x"0F5D1",
									 x"0FF18",x"0FFBE",x"0FFDF",x"0FFFF",x"10022",x"0FFFF",x"10022",x"0FFDF",x"0FF9D",x"0FF1A",
									 x"0EE34",x"0ECCB",x"0E425",x"0EC03",x"0F421",x"0F462",x"0F4A3",x"0F4C4",x"0FCE4",x"0FD04",
									 x"0FD25",x"0FD45",x"0FD64",x"0FD84",x"0FD85",x"0FDA5",x"10000",x"0FDC5",x"10000",x"0FDE8",
									 x"0FE4B",x"0FED0",x"0FF34",x"0FF56",x"0FF36",x"10000",x"0FF35",x"0FF56",x"10002",x"0FF36",
									 x"0FF56",x"10000",x"0FF36",x"10001",x"0FF56",x"10008",x"0FF36",x"10000",x"0FF56",x"1004E",
									 x"0FF36",x"10000",x"0FF56",x"10008",x"0FF36",x"10003",x"0FF56",x"10000",x"0FF36",x"10001",
									 x"0FF56",x"0FF55",x"10000",x"0FF76",x"0FF56",x"0FF15",x"0FEB0",x"0FE4B",x"0FE07",x"0FDC6",
									 x"0FD85",x"0FDA5",x"10001",x"0FD65",x"0FD64",x"0FD44",x"0FD24",x"10000",x"0FD04",x"0F4C3",
									 x"0FCA3",x"0F463",x"0F423",x"0F403",x"0F425",x"0ECAA",x"0F5F2",x"0FEF9",x"0FF9D",x"0FFDF",
									 x"0FFFF",x"10021",x"0FFFF",x"10022",x"0FFBE",x"0FF1A",x"0F654",x"0ED2C",x"0EC66",x"0EC24",
									 x"0F443",x"0F462",x"0F4A2",x"0F4E3",x"0F4E4",x"0FD04",x"0FD24",x"0FD44",x"0FD64",x"0FD65",
									 x"0F585",x"0FDA5",x"10000",x"0FDC4",x"0FDC5",x"0FDE7",x"0FE4C",x"0FEB0",x"0FF13",x"0FF56",
									 x"0FF36",x"10007",x"0FF35",x"10001",x"0FF56",x"1000A",x"0FF36",x"10003",x"0FF56",x"10005",
									 x"0FF36",x"10036",x"0FF56",x"1000C",x"0FF36",x"10002",x"0FF56",x"10000",x"0FF36",x"1000D",
									 x"0FF56",x"0FF36",x"10000",x"0FF35",x"0FF55",x"0FF56",x"0FF36",x"0FF14",x"0FEB0",x"0FE6C",
									 x"0FDE9",x"0FD85",x"0FD84",x"0FDA5",x"10000",x"0FD84",x"0FD64",x"10000",x"0FD44",x"0FD24",
									 x"0FD04",x"0FCE3",x"0F4C3",x"10000",x"0F483",x"0F443",x"0F403",x"0EC26",x"0ED0C",x"0F613",
									 x"0FEF9",x"0FF9D",x"0F7DF",x"0FFFF",x"10020",x"0FFFF",x"10022",x"0FF7C",x"0F695",x"0F56E",
									 x"0EC68",x"0EC24",x"0F423",x"0FC63",x"0FCA3",x"0F4C3",x"0F4E3",x"0FD04",x"0FD24",x"0FD45",
									 x"0FD65",x"0FD85",x"10001",x"0FDA5",x"0FDC4",x"10000",x"0FE07",x"0FE2B",x"0FEB0",x"0FF13",
									 x"0FF35",x"0FF56",x"10000",x"0FF35",x"0FF36",x"10004",x"0FF35",x"10002",x"0FF55",x"0FF56",
									 x"10009",x"0FF36",x"10003",x"0FF56",x"10005",x"0FF36",x"10031",x"0FF56",x"0FF55",x"10002",
									 x"0FF56",x"1000C",x"0FF36",x"10002",x"0FF56",x"10004",x"0FF36",x"10000",x"0FF55",x"10003",
									 x"0FF56",x"0FF36",x"10004",x"0FF35",x"10000",x"0FF36",x"10000",x"0FF35",x"0FF13",x"0FED1",
									 x"0FE4C",x"0FDE7",x"0FDC4",x"0FDA4",x"0FDA5",x"10000",x"0FD85",x"0FD64",x"0FD44",x"10000",
									 x"0FD24",x"0FD04",x"10000",x"0F4E4",x"0F4A3",x"0F463",x"0F423",x"0EC23",x"0EC87",x"0F54E",
									 x"0FE34",x"0FF3A",x"0FFFF",x"0F7FF",x"0FFFF",x"1001F",x"0FFFF",x"10021",x"0FFBD",x"0F6D6",
									 x"0ED8F",x"0F488",x"0F404",x"0F442",x"10000",x"0FC83",x"0FCC3",x"0FD04",x"0F504",x"0FD24",
									 x"0FD44",x"0FD65",x"0FD85",x"10000",x"0FDA5",x"0FD85",x"0FDA4",x"0FDC4",x"0FE06",x"0FE49",
									 x"0FE8F",x"0FEF3",x"0FF35",x"0FF56",x"10000",x"0FF36",x"0FF35",x"10009",x"0FF55",x"0FF56",
									 x"0FF55",x"10064",x"0FF35",x"0FF55",x"10002",x"0FF35",x"10001",x"0FF55",x"10001",x"0FF35",
									 x"10004",x"0FF36",x"10000",x"0FF55",x"0FF15",x"0FEB0",x"0F64A",x"0FE06",x"0FDC5",x"0FDA5",
									 x"10001",x"0FD85",x"0FD65",x"10000",x"0FD44",x"0FD24",x"0F504",x"0F4E4",x"0F4C3",x"0F483",
									 x"0F443",x"0F422",x"0F424",x"0F488",x"0F52E",x"0FE96",x"0FFBD",x"0F7DE",x"0FFFF",x"1001F",
									 x"0FFFF",x"1001F",x"0FFDF",x"0FF9D",x"0FEF8",x"0F5D0",x"0ECA8",x"0F424",x"0F422",x"0F462",
									 x"0F483",x"0F4A3",x"0FCE4",x"0FD24",x"0F524",x"0FD44",x"10000",x"0FD85",x"10000",x"0FDA5",
									 x"10000",x"0FDA4",x"0FDA5",x"0FDE7",x"0FE49",x"0FE8D",x"0FEF2",x"0FF35",x"0FF56",x"0FF36",
									 x"0FF35",x"1000A",x"0FF55",x"10067",x"0FF35",x"1000F",x"0FF16",x"0FF36",x"0FF56",x"0FF36",
									 x"0FEF3",x"0FE8E",x"0FE4A",x"0FE07",x"0FDC6",x"0FDA5",x"10001",x"0FD85",x"0FD65",x"0FD45",
									 x"0FD44",x"0F524",x"0F504",x"0FD04",x"0FCC4",x"0F483",x"0FC62",x"0F422",x"0F424",x"0F468",
									 x"0F5AF",x"0FEF8",x"0FF9C",x"0FFFF",x"1001F",x"0FFFF",x"1001F",x"0FFBE",x"0FEF9",x"0FE13",
									 x"0F4EB",x"0EC25",x"0F423",x"0F463",x"0F483",x"0F4A3",x"0F4C4",x"0F504",x"0F524",x"10000",
									 x"0FD44",x"0FD65",x"0FD85",x"0FDA5",x"0FDC5",x"10001",x"0FDC7",x"0FE0A",x"0FE8D",x"0FEF1",
									 x"0FF34",x"0FF36",x"0FF16",x"0FF15",x"0FF35",x"10000",x"0FF15",x"10002",x"0FF35",x"10004",
									 x"0FF55",x"10010",x"0FF35",x"10005",x"0FF55",x"10000",x"0FF35",x"10020",x"0FF55",x"10001",
									 x"0FF35",x"10007",x"0FF55",x"10002",x"0FF35",x"10003",x"0FF55",x"10005",x"0FF35",x"10006",
									 x"0FF55",x"10007",x"0FF35",x"1000C",x"0FF34",x"10000",x"0FF15",x"10000",x"0FF34",x"0FF15",
									 x"0FF35",x"0FED2",x"0FE8F",x"0FE2B",x"0FDC7",x"0FDC5",x"10000",x"0FDA5",x"10000",x"0FD85",
									 x"0FD65",x"0FD64",x"10000",x"0F524",x"0F504",x"0FCE3",x"0FCA3",x"0F483",x"0F442",x"0F422",
									 x"0F424",x"0F4CA",x"0FDF2",x"0FEF9",x"0FF9D",x"0FFFF",x"1001E",x"0FFFF",x"1001D",x"0FFDF",
									 x"0FFDE",x"0FF7C",x"0F675",x"0F54E",x"0F447",x"0F403",x"0F443",x"0EC83",x"0F4A3",x"0F4C4",
									 x"0F4E4",x"0F504",x"0FD24",x"0FD44",x"0FD64",x"0FD85",x"0FDA5",x"0FDC5",x"10000",x"0FDE5",
									 x"0FDC5",x"0FDE8",x"0FE6D",x"0FED1",x"0FF13",x"0FF35",x"0FF16",x"0FF15",x"10000",x"0FF14",
									 x"10000",x"0FF15",x"0FF14",x"10001",x"0FF34",x"0FF35",x"10003",x"0FF55",x"1000B",x"0FF34",
									 x"0FF35",x"10001",x"0FF34",x"0FF55",x"10004",x"0FF35",x"0FF34",x"10000",x"0FF35",x"0FF55",
									 x"1001F",x"0FF35",x"10001",x"0FF55",x"10017",x"0FF35",x"10004",x"0FF55",x"10008",x"0FF35",
									 x"1000A",x"0FF34",x"0FF35",x"10000",x"0FF34",x"10000",x"0FF15",x"10000",x"0FF34",x"0FF14",
									 x"0FF35",x"0FEF4",x"0FED2",x"0FE6D",x"0FDE8",x"0FDC6",x"0FDC5",x"10000",x"0FDA5",x"10000",
									 x"0FD85",x"0FD65",x"0FD64",x"0FD44",x"0F524",x"0FCE4",x"0FCC3",x"0F4A4",x"0F483",x"0F442",
									 x"0F402",x"0EC46",x"0F50D",x"0F635",x"0FF3B",x"0FFBE",x"0FFFF",x"1001D",x"0FFFF",x"1001C",
									 x"0FFDE",x"0FFDF",x"0FF9C",x"0EEB6",x"0ED6F",x"0EC89",x"0F404",x"0F422",x"0F463",x"0F4A3",
									 x"0F4E4",x"0FD04",x"10000",x"0FD24",x"0FD44",x"0FD64",x"10000",x"0FD86",x"0FDA6",x"0FDC5",
									 x"10001",x"0FDE6",x"0FE2B",x"0FED0",x"0FF13",x"0FF35",x"0FF15",x"10002",x"0FF14",x"0FF34",
									 x"10007",x"0FF54",x"10003",x"0FF34",x"1000B",x"0FF54",x"10003",x"0FF34",x"10011",x"0FF54",
									 x"10009",x"0FF34",x"10006",x"0FF54",x"10003",x"0FF34",x"10005",x"0FF54",x"1000F",x"0FF34",
									 x"10005",x"0FF54",x"10009",x"0FF34",x"1000E",x"0FF35",x"10000",x"0FF15",x"10000",x"0FF34",
									 x"0FF15",x"0FF14",x"0FED0",x"0FE4B",x"0FDE7",x"0FDC6",x"0FDA5",x"0FDC5",x"0FDA5",x"0FDA6",
									 x"0FD85",x"0FD64",x"0FD44",x"0FD24",x"10000",x"0F504",x"0F4C4",x"0F4A3",x"0F462",x"0F422",
									 x"0EC23",x"0EC66",x"0ED4D",x"0F675",x"0FF5C",x"0FFDE",x"0FFFF",x"1001C",x"0FFFF",x"1001C",
									 x"0FFDF",x"0FF9E",x"0FF19",x"0E5D1",x"0E4C9",x"0EC25",x"0F402",x"0F461",x"0F4A2",x"0F4C3",
									 x"0F4E4",x"0FD04",x"0FD24",x"0FD45",x"0FD65",x"0FD85",x"10000",x"0FDA6",x"10000",x"0FDC5",
									 x"10000",x"0FDE6",x"0FE29",x"0FE6D",x"0FEF2",x"0FF34",x"10000",x"0FF35",x"0FF15",x"10000",
									 x"0FF14",x"0FF34",x"10085",x"0FF15",x"10000",x"0FF14",x"0FF34",x"0FF35",x"0FF15",x"0FEF2",
									 x"0FEAE",x"0FE49",x"0FDE7",x"0FDC5",x"0FDA5",x"10000",x"0FDA6",x"0FDA5",x"0FD85",x"0FD64",
									 x"0FD44",x"0FD24",x"0FD04",x"0F504",x"0F4C3",x"0F482",x"0FC62",x"0EC22",x"0EC23",x"0ECA8",
									 x"0F590",x"0FED9",x"0F79D",x"0FFFF",x"1001C",x"0FFFF",x"1001A",x"0FFDF",x"0FFFF",x"0FFBF",
									 x"0FF3B",x"0FE54",x"0ED2C",x"0EC66",x"0F424",x"0F422",x"0F482",x"0F4C3",x"0F4E4",x"0F504",
									 x"0FD24",x"10000",x"0FD44",x"0FD85",x"10000",x"0FDA5",x"0FDC6",x"10000",x"0FDC5",x"0FDE6",
									 x"0FE29",x"0FE6D",x"0FED1",x"0FF14",x"0FF34",x"10002",x"0FF14",x"0FF34",x"10087",x"0FF14",
									 x"0FF34",x"10001",x"0FF35",x"0FF34",x"0FEF1",x"0FE8C",x"0FE29",x"0FDE6",x"0FDC5",x"10001",
									 x"0FDA5",x"10000",x"0FD65",x"10000",x"0FD44",x"0FD24",x"0F524",x"0F4E4",x"0F4A3",x"0FC83",
									 x"0F442",x"0EC22",x"0F445",x"0F4EB",x"0FE55",x"0FF1A",x"0FFBD",x"0FFFF",x"1001B",x"0FFFF",
									 x"1001C",x"0FF7C",x"0FE76",x"0F56E",x"0EC87",x"0EC24",x"0FC44",x"0F463",x"0F4A3",x"0F4E4",
									 x"10000",x"0F524",x"0FD44",x"10000",x"0FD64",x"0FD85",x"0FDA5",x"0FDC5",x"0FDC6",x"10000",
									 x"0FDE6",x"0F608",x"0FE6C",x"0FED0",x"0FEF3",x"0FF15",x"0FF34",x"10000",x"0FF14",x"10000",
									 x"0FF34",x"1002E",x"0FF14",x"10003",x"0FF34",x"10054",x"0FF14",x"0FF33",x"0FF34",x"0FF35",
									 x"10000",x"0FF13",x"0FED0",x"0FE6C",x"0FE28",x"0FDE6",x"0FDC5",x"0FDC6",x"0FDC5",x"0FDA5",
									 x"0FD85",x"0FD65",x"10000",x"0FD45",x"0F525",x"0F504",x"0F4C4",x"0F4A3",x"0F463",x"0F443",
									 x"0F423",x"0EC67",x"0F54E",x"0FE55",x"0FF5A",x"0FFDE",x"0FFFF",x"1001A",x"0FFFF",x"1001A",
									 x"0FFDF",x"0FFBC",x"0F6D7",x"0F5B0",x"0EC88",x"0EC23",x"0EC22",x"0FC63",x"0FCA3",x"0F4E3",
									 x"0F504",x"0FD04",x"0FD44",x"0FD64",x"0FD85",x"10000",x"0FDA5",x"0FDC5",x"10000",x"0FDC6",
									 x"0FDE6",x"0FE07",x"0FE4B",x"0FED0",x"0FF12",x"0FF14",x"0FF15",x"0FF13",x"10002",x"0FF33",
									 x"10000",x"0FF34",x"10002",x"0FF33",x"10006",x"0FF34",x"10010",x"0FF33",x"10001",x"0FF34",
									 x"10011",x"0FF33",x"10009",x"0FF34",x"10006",x"0FF33",x"10002",x"0FF34",x"10006",x"0FF33",
									 x"1000F",x"0FF34",x"10005",x"0FF33",x"10007",x"0FF34",x"1000A",x"0FF33",x"10000",x"0FF34",
									 x"10005",x"0FF14",x"0FF33",x"0FF13",x"0FF14",x"10001",x"0FF13",x"0FECF",x"0FE6B",x"0FE07",
									 x"0FE06",x"0FDC6",x"0FDC5",x"10000",x"0FDA5",x"0FD85",x"0FD65",x"10000",x"0FD44",x"0FD24",
									 x"0FD04",x"0FCC3",x"0F4A3",x"0F463",x"0EC42",x"0EC44",x"0EC88",x"0F56E",x"0FE96",x"0FF9D",
									 x"0FFDF",x"0FFFF",x"10019",x"0FFFF",x"10019",x"0FFDF",x"0FFFF",x"0FF7B",x"0F612",x"0F52C",
									 x"0EC45",x"0F442",x"0EC42",x"0F483",x"0F4C3",x"0F503",x"0FD03",x"0FD24",x"0FD64",x"0FD85",
									 x"10000",x"0FDA5",x"10001",x"0FDC5",x"10000",x"0FDE6",x"0FE28",x"0FE8D",x"0FEF2",x"0FF13",
									 x"0FF14",x"10001",x"0FF13",x"10001",x"0FF33",x"10000",x"0FF34",x"10001",x"0FF33",x"0FF13",
									 x"1000A",x"0FF14",x"10009",x"0FF13",x"10004",x"0FF14",x"0FF34",x"10001",x"0FF14",x"1000C",
									 x"0FF13",x"1000B",x"0FF14",x"10004",x"0FF13",x"10004",x"0FF14",x"10004",x"0FF13",x"10011",
									 x"0FF14",x"10003",x"0FF13",x"1000B",x"0FF14",x"10003",x"0FF13",x"0FF33",x"10004",x"0FF34",
									 x"10001",x"0FF14",x"0FF13",x"10000",x"0FF14",x"0FF13",x"10000",x"0FF14",x"10002",x"0FF11",
									 x"0FEAC",x"0FE49",x"0FE07",x"0FDC6",x"0FDC5",x"10000",x"0FDA5",x"0FD85",x"10000",x"0FD65",
									 x"0FD43",x"10000",x"0FD23",x"0FCE3",x"0F4C3",x"0F482",x"0EC82",x"0EC43",x"0EC25",x"0F4EA",
									 x"0F5F2",x"0F73B",x"0FFDF",x"10000",x"0FFFF",x"10018",x"0FFFF",x"10019",x"0FFDF",x"0FF9D",
									 x"0FED6",x"0F56E",x"0EC88",x"0EC24",x"0EC42",x"0F483",x"0F4A3",x"0F4E3",x"0F504",x"0FD24",
									 x"0FD44",x"0FD64",x"0FD85",x"10000",x"0FDA5",x"0FDC5",x"10002",x"0FE07",x"0F64A",x"0FEAF",
									 x"0FEF2",x"0FF14",x"0FEF4",x"0FF13",x"10093",x"0FF14",x"10000",x"0FEF3",x"0FECF",x"0FE8B",
									 x"0FE28",x"0FDE6",x"0FDC5",x"0FDA5",x"0FDC5",x"0FDA5",x"0FD85",x"10000",x"0FD65",x"0FD44",
									 x"0FD24",x"10000",x"0FCE4",x"0F4A3",x"0F483",x"0F443",x"0EC23",x"0EC66",x"0ED2D",x"0F697",
									 x"0FF7D",x"0FFDF",x"0FFFF",x"10018",x"0FFFF",x"10018",x"0FFDF",x"0FFBE",x"0FF1A",x"0F5F1",
									 x"0EC88",x"0F424",x"0F422",x"0F462",x"0F4A3",x"0FCE3",x"0FD04",x"0FD24",x"0FD44",x"0FD64",
									 x"0FD85",x"10000",x"0FDA5",x"10000",x"0FDC6",x"10001",x"0FDE7",x"0FE4A",x"0FE8D",x"0FED1",
									 x"0FEF3",x"0FF13",x"0FEF3",x"10000",x"0FF13",x"10095",x"0FEF1",x"0FEAE",x"0FE6A",x"0FE07",
									 x"0FDC5",x"10002",x"0FDA5",x"0FD85",x"10000",x"0FD65",x"0FD44",x"0FD24",x"0FD04",x"0FCC3",
									 x"10000",x"0F482",x"0EC42",x"0EC23",x"0E488",x"0EDD0",x"0F719",x"0F7BD",x"0FFFF",x"0FFFE",
									 x"10000",x"0FFFF",x"10015",x"0FFFF",x"10018",x"0FFDE",x"0FF7C",x"0F697",x"0ED4D",x"0F424",
									 x"0FC02",x"0FC42",x"0F483",x"0F4C3",x"0F4E3",x"0FD04",x"0FD24",x"0FD64",x"0FD65",x"0FD85",
									 x"0FDA5",x"10000",x"0FDC6",x"0FDE6",x"10000",x"0FDE7",x"0FE29",x"0FE8C",x"0FED0",x"0FEF2",
									 x"0FF14",x"0FEF3",x"10002",x"0FF13",x"10091",x"0FEF3",x"0FF13",x"10000",x"0FEF3",x"0FED1",
									 x"0FE8D",x"0FE49",x"0FDE6",x"0FDC5",x"10001",x"0FDA6",x"0FD86",x"0FD85",x"0FD65",x"0FD45",
									 x"0FD44",x"0FD04",x"0FCE3",x"0FCC3",x"0F4A2",x"0F462",x"0EC22",x"0EC45",x"0ED2B",x"0F695",
									 x"0F77B",x"0F7DE",x"10000",x"0FFFE",x"0FFFF",x"10015",x"0FFFF",x"10016",x"0F7FF",x"0FFFE",
									 x"0FF7C",x"0FEF9",x"0EDF3",x"0E4C9",x"0EC23",x"0F422",x"0F463",x"0F4C4",x"0F4E3",x"0FD04",
									 x"0FD24",x"0FD44",x"0FD84",x"0FD85",x"0FDA5",x"0FDC5",x"10000",x"0FDC6",x"0FDE6",x"10000",
									 x"0FE08",x"0FE4B",x"0FEAF",x"0FED2",x"0FEF3",x"10000",x"0FEF2",x"10002",x"0FEF3",x"10000",
									 x"0FEF2",x"10001",x"0FF13",x"10086",x"0FF12",x"10002",x"0FEF2",x"10002",x"0FEF3",x"0FF14",
									 x"0FEF3",x"0FEAF",x"0FE6B",x"0FE08",x"0FDE6",x"10000",x"0FDC5",x"10000",x"0FDA6",x"0FDA5",
									 x"0FD85",x"0FD64",x"0FD44",x"0FD24",x"0F503",x"0FCE3",x"0F4A3",x"0F463",x"0F422",x"0EC24",
									 x"0EC87",x"0F5D0",x"0F6D8",x"0F77D",x"0F7BF",x"0FFFF",x"10016",x"0FFFF",x"10016",x"0F7DF",
									 x"0FFBD",x"0FF19",x"0FE55",x"0ED4E",x"0E466",x"0EC22",x"0F442",x"0F483",x"0F4C4",x"0F4E3",
									 x"0FD24",x"0FD44",x"0FD64",x"0FD85",x"0FDA5",x"10000",x"0FDC6",x"10000",x"0FDE6",x"10000",
									 x"0FE06",x"0FE29",x"0FE6D",x"0FED1",x"0FEF3",x"10000",x"0FEF2",x"10008",x"0FF12",x"10089",
									 x"0FEF2",x"10003",x"0FEF3",x"0FF13",x"10000",x"0FED1",x"0FE8E",x"0FE29",x"0FDE7",x"0FDE6",
									 x"0FDC5",x"10001",x"0FDA5",x"10000",x"0FD85",x"0FD64",x"0FD44",x"0FD24",x"0FD04",x"0F4C4",
									 x"0F4A3",x"0FC63",x"0F443",x"0EC24",x"0F50B",x"0F613",x"0F6FA",x"0FFBE",x"0FFDF",x"10000",
									 x"0FFFF",x"10014",x"0FFFF",x"10014",x"0FFDE",x"0F7DF",x"10000",x"0FF9C",x"0F675",x"0ED4F",
									 x"0EC88",x"0EC44",x"0F462",x"10000",x"0F4A3",x"0F504",x"0F503",x"0FD24",x"0FD44",x"0FD84",
									 x"0FDA5",x"10001",x"0FDC6",x"10001",x"0FDE6",x"0FE27",x"0FE4A",x"0FEAE",x"0FED2",x"0FEF3",
									 x"0FEF2",x"0FEF1",x"10000",x"0FEF2",x"1000A",x"0FF12",x"1007C",x"0FEF2",x"10005",x"0FF11",
									 x"0FF12",x"10000",x"0FEF2",x"10005",x"0FEF1",x"0FEB0",x"0FE6B",x"0FE08",x"0FDE6",x"0FDE5",
									 x"10001",x"0FDC5",x"0FDA5",x"10000",x"0FD85",x"0FD64",x"0FD44",x"0FD23",x"0F4E3",x"0F4C3",
									 x"0FC82",x"0F462",x"0EC23",x"0EC67",x"0ED2D",x"0EE55",x"0FF7C",x"0FFBE",x"0FFDE",x"0FFDF",
									 x"0FFFF",x"10013",x"0FFFF",x"10014",x"0FFDF",x"0F7DF",x"0F7BE",x"0FF5B",x"0EDD1",x"0EC89",
									 x"0F445",x"0F423",x"0F463",x"0F4A3",x"0F4E3",x"0F504",x"0F524",x"0FD44",x"0FD64",x"0FD85",
									 x"10000",x"0FDA5",x"0FDC6",x"10000",x"0FDC5",x"0FDE6",x"0FE07",x"0FE28",x"0FE6C",x"0FED0",
									 x"0FEF3",x"10000",x"0FEF2",x"10000",x"0FEF1",x"10001",x"0FEF2",x"10019",x"0FF12",x"10023",
									 x"0FEF2",x"10004",x"0FF12",x"1001D",x"0FEF2",x"10009",x"0FF12",x"1000B",x"0FEF2",x"10014",
									 x"0FEF1",x"10000",x"0FEF2",x"10002",x"0FEF1",x"0FED1",x"0FE8D",x"0FE2A",x"0FE07",x"0FDE5",
									 x"10001",x"0FDC5",x"10000",x"0FDA5",x"10000",x"0FD84",x"0F564",x"0FD24",x"0F504",x"0F4C3",
									 x"0F4A3",x"0F463",x"0F442",x"0EC44",x"0EC68",x"0F5B0",x"0F719",x"0F7BE",x"0F7DE",x"0FFDF",
									 x"0FFFF",x"10013",x"0FFFF",x"10015",x"0FFDF",x"0FF9E",x"0FED8",x"0ED4D",x"0EC45",x"0EC23",
									 x"0F443",x"0FC83",x"0F4A2",x"0F4E3",x"0F524",x"0FD44",x"0FD64",x"0FD65",x"0FD85",x"0FDA5",
									 x"10000",x"0FDC6",x"0FDE6",x"0FDE5",x"0FE06",x"0FE28",x"0FE4A",x"0FE8E",x"0FED1",x"0FEF3",
									 x"0FEF2",x"0FEF1",x"10006",x"0FEF2",x"1001F",x"0FF12",x"10002",x"0FEF2",x"10012",x"0FF12",
									 x"10002",x"0FEF2",x"1001C",x"0FF12",x"10002",x"0FEF2",x"1000C",x"0FF12",x"10008",x"0FEF2",
									 x"10013",x"0FEF1",x"10007",x"0FEF2",x"10000",x"0FED1",x"0FEAE",x"0FE4B",x"0FE27",x"0FE05",
									 x"0FDE5",x"0FDE6",x"0FDC6",x"0FDC5",x"10000",x"0FDA5",x"0FD84",x"0FD64",x"0FD44",x"0FD04",
									 x"0FCE4",x"0F4C3",x"0F483",x"0F462",x"0F443",x"0EC45",x"0ED4C",x"0F6B6",x"0FF9C",x"0FFDE",
									 x"10000",x"0FFFF",x"10013",x"0FFFF",x"10014",x"0F7FF",x"0FFBE",x"0FF1B",x"0F613",x"0ECA8",
									 x"0F423",x"0EC42",x"0F482",x"0FCA3",x"0FCE3",x"0F504",x"0F524",x"0FD44",x"0FD85",x"10000",
									 x"0FDA5",x"0FDC5",x"0FDC6",x"10000",x"0FDE6",x"10000",x"0FE07",x"0FE29",x"0FE6C",x"0FEAF",
									 x"0FED2",x"0FED3",x"0FEF2",x"0FEF1",x"1009C",x"0FEF2",x"10000",x"0FEB0",x"0FE6C",x"0FE48",
									 x"0FE06",x"0FDE6",x"0FDE7",x"0FDC6",x"0FDC5",x"10000",x"0FDA5",x"10000",x"0FD84",x"0FD44",
									 x"0FD24",x"0FD04",x"0FCE3",x"0F4A3",x"0F483",x"0F442",x"0EC22",x"0EC87",x"0EDB0",x"0FF1A",
									 x"0FF9D",x"0FFDE",x"0FFFF",x"10013",x"0FFFF",x"10013",x"0F7FF",x"0F7DF",x"0FF3B",x"0FE97",
									 x"0ED2E",x"0EC44",x"0F421",x"0F462",x"0FCA3",x"0FCC3",x"0FD03",x"0FD24",x"0FD44",x"0FD64",
									 x"0FD85",x"0FDA5",x"10000",x"0FDC6",x"0FDE6",x"10000",x"0FE05",x"0FE06",x"0FE28",x"0FE4A",
									 x"0FE8E",x"0FED0",x"0FED2",x"10000",x"0FED1",x"0FEF0",x"0FEF1",x"1009A",x"0FED1",x"0FEF2",
									 x"0FED1",x"10000",x"0FEAE",x"0FE6A",x"0FE27",x"0FDE6",x"0FDC6",x"10002",x"0FDC5",x"0FDA5",
									 x"0FD85",x"0FD64",x"0FD44",x"0FD24",x"0FD04",x"0FCC3",x"0F4A3",x"0F463",x"0F402",x"0EC25",
									 x"0ECEC",x"0F656",x"0FF1B",x"0FFBE",x"0FFDF",x"0FFFF",x"10012",x"0FFFF",x"10012",x"0FFDF",
									 x"10000",x"0FFBE",x"0FED8",x"0FE33",x"0ECCA",x"0EC03",x"0FC42",x"0F483",x"0FCC3",x"0FCE4",
									 x"0FD04",x"0FD24",x"0FD64",x"0FD85",x"10000",x"0FDA5",x"0FDC5",x"0FDC6",x"0FDE6",x"10000",
									 x"0FE05",x"0FE26",x"0FE48",x"0FE6C",x"0FEAF",x"0FED0",x"0FED1",x"10000",x"0FED0",x"0FEF0",
									 x"0FEF1",x"1000B",x"0FF11",x"10001",x"0FEF1",x"10011",x"0FF11",x"10001",x"0FEF1",x"10007",
									 x"0FF11",x"10000",x"0FEF1",x"10008",x"0FF11",x"10001",x"0FEF1",x"10002",x"0FF11",x"0FEF1",
									 x"10030",x"0FF11",x"10006",x"0FEF1",x"1001D",x"0FED1",x"10002",x"0FECF",x"0FE8C",x"0FE49",
									 x"0FE07",x"0FDE6",x"10002",x"0FDC6",x"0FDA5",x"0FD85",x"10000",x"0FD64",x"0FD24",x"0FD04",
									 x"0FCE3",x"0FCC3",x"0F483",x"0F422",x"0F403",x"0EC89",x"0F5F2",x"0FEB8",x"0FF9D",x"0FFDF",
									 x"10000",x"0FFFF",x"10011",x"0FFFF",x"10011",x"0FFDF",x"0F7BE",x"0FFDF",x"0FF7D",x"0F634",
									 x"0F58E",x"0E467",x"0EC23",x"0F442",x"0F483",x"0FCC4",x"0FCE4",x"0FD24",x"0FD44",x"0FD64",
									 x"0FD85",x"0FDA5",x"10000",x"0FDC6",x"0FDE6",x"10000",x"0FE06",x"0FE05",x"0FE26",x"0FE49",
									 x"0FE8D",x"0FED0",x"0FEF0",x"0FEF1",x"0FED0",x"10000",x"0FEF0",x"0FEF1",x"10006",x"0FEF0",
									 x"10000",x"0FEF1",x"10001",x"0FEF0",x"10017",x"0FEF1",x"10001",x"0FEF0",x"10019",x"0FEF1",
									 x"10000",x"0FEF0",x"1002B",x"0FEF1",x"0FEF0",x"1001C",x"0FEF1",x"10002",x"0FEF0",x"10000",
									 x"0FEF1",x"0FED1",x"10002",x"0FED0",x"10000",x"0FEF0",x"0FED0",x"0FE8E",x"0FE4B",x"0FE08",
									 x"0FE05",x"0FDE6",x"10001",x"0FDC6",x"0FDA6",x"0FDA5",x"0FD85",x"0FD84",x"0FD44",x"0FD24",
									 x"0FD04",x"0FCC3",x"0F483",x"0F462",x"0F422",x"0EC65",x"0ED4D",x"0EE33",x"0FF7C",x"0FFDF",
									 x"10000",x"0FFFF",x"10011",x"0FFFF",x"10011",x"0FFDE",x"0F7DE",x"0F7BF",x"0FF1B",x"0ED8F",
									 x"0ECC7",x"0EC64",x"0F442",x"0FC82",x"0FCA3",x"0FCC4",x"0FD04",x"0FD44",x"0F544",x"0FD85",
									 x"10000",x"0FDA5",x"10000",x"0FDC5",x"0FDE6",x"10000",x"0FE06",x"0FE05",x"0FE27",x"0FE6B",
									 x"0FEAF",x"0FED0",x"0FEF0",x"0FED0",x"10001",x"0FEF0",x"1009C",x"0FED0",x"10002",x"0FEAF",
									 x"0FE6C",x"0FE28",x"0FE05",x"0FDE6",x"10001",x"0FDC5",x"0FDA5",x"10000",x"0FD85",x"0FD65",
									 x"0FD64",x"0FD44",x"0FD24",x"0FCE3",x"0FCA3",x"0FC83",x"0F442",x"0F443",x"0ECA8",x"0ED4E",
									 x"0FEF8",x"0FFBE",x"0F7DF",x"0FFDF",x"0FFFF",x"10010",x"0FFFF",x"10011",x"0FFDF",x"0FFBE",
									 x"0FF7D",x"0F697",x"0ECEB",x"0EC25",x"0F424",x"0FC63",x"0FC82",x"0FCA3",x"0FCE4",x"0FD24",
									 x"0FD44",x"0FD64",x"0FD85",x"10000",x"0FDA5",x"10000",x"0FDC6",x"0FDE6",x"10000",x"0FDE5",
									 x"0FE05",x"0FE28",x"0FE8C",x"0FEAF",x"0FED0",x"10003",x"0FEF0",x"0FED0",x"10000",x"0FEF0",
									 x"10006",x"0FED0",x"10004",x"0FEF0",x"10010",x"0FED0",x"10005",x"0FEF0",x"10003",x"0FED0",
									 x"10005",x"0FEF0",x"10000",x"0FED0",x"1000E",x"0FEF0",x"1000D",x"0FED0",x"10004",x"0FEF0",
									 x"10016",x"0FED0",x"10011",x"0FEF0",x"1000D",x"0FED0",x"10004",x"0FEF0",x"0FED0",x"10002",
									 x"0FEAF",x"0FE8D",x"0FE29",x"0FE06",x"10001",x"0FDE6",x"0FDC6",x"10000",x"0FDA5",x"0FD85",
									 x"10000",x"0FD64",x"10000",x"0FD44",x"0FD04",x"0FCC3",x"0FC83",x"0F442",x"0F423",x"0E446",
									 x"0ECCB",x"0F676",x"0F77C",x"0F7DF",x"0FFDF",x"0FFFF",x"10010",x"0FFFF",x"10010",x"0FFDF",
									 x"10000",x"0FF9E",x"0FF1B",x"0F613",x"0EC88",x"0F3E3",x"0FC23",x"0FC63",x"0FCA3",x"0FCC3",
									 x"0FD04",x"0FD24",x"0FD64",x"0FD65",x"0FD85",x"0FDA5",x"10000",x"0FDC6",x"0FDE6",x"10001",
									 x"0FDE5",x"0FE06",x"0FE49",x"0FE8D",x"0FED0",x"100A7",x"0FEAE",x"0FE4A",x"0FE27",x"0FE06",
									 x"10001",x"0FDE6",x"0FDC6",x"0FDC5",x"0FDA5",x"0FD85",x"10000",x"0FD64",x"0FD44",x"0FD04",
									 x"0FCE3",x"0FCA3",x"0FC83",x"0F443",x"0EC24",x"0EC68",x"0F5B2",x"0F71A",x"0F79E",x"0F7DF",
									 x"0FFFF",x"10010",x"0FFFF",x"10010",x"0FFDF",x"0FFBE",x"0FF5C",x"0F6B7",x"0E54D",x"0EC66",
									 x"0F403",x"0F443",x"0F484",x"0F4E3",x"0FCE3",x"0FD24",x"0FD44",x"0FD64",x"0FD85",x"0FDA5",
									 x"10000",x"0FDC5",x"0FDC6",x"0FDE6",x"0FE06",x"10000",x"0FE26",x"0FE27",x"0FE6A",x"0FEAF",
									 x"0FED1",x"0FED0",x"10045",x"0FEF0",x"10000",x"0FED0",x"10015",x"0FEF0",x"10000",x"0FED0",
									 x"10043",x"0FEF1",x"0FECF",x"0FE6B",x"0FE48",x"0FE27",x"0FE06",x"10001",x"0FDE6",x"0FDC6",
									 x"0FDA5",x"10000",x"0FD85",x"10000",x"0FD44",x"0FD24",x"0FCE3",x"0FCC3",x"0FC83",x"0FC63",
									 x"0F423",x"0EC05",x"0ED0D",x"0F676",x"0FF5C",x"0F7BF",x"0FFDF",x"0FFFF",x"1000F",x"0FFFF",
									 x"10010",x"0FFDF",x"0FF9D",x"0FF3A",x"0F634",x"0E4A9",x"0EC44",x"0EC22",x"0EC63",x"0F4A4",
									 x"0F4E3",x"0F503",x"0FD24",x"0FD64",x"10000",x"0FD85",x"0FDA5",x"10000",x"0FDC5",x"0FDE6",
									 x"10000",x"0FE06",x"10001",x"0FE48",x"0FE8C",x"0FECF",x"0FED0",x"0FECF",x"10000",x"0FED0",
									 x"10000",x"0FECF",x"10001",x"0FED0",x"1000A",x"0FECF",x"10005",x"0FED0",x"0FECF",x"0FED0",
									 x"1000A",x"0FECF",x"10002",x"0FED0",x"10001",x"0FECF",x"10001",x"0FED0",x"10001",x"0FECF",
									 x"10000",x"0FED0",x"10008",x"0FECF",x"10008",x"0FED0",x"10012",x"0FECF",x"10001",x"0FED0",
									 x"10010",x"0FECF",x"0FED0",x"10004",x"0FECF",x"10001",x"0FED0",x"10000",x"0FECF",x"10008",
									 x"0FED0",x"10010",x"0FECF",x"10008",x"0FED0",x"10000",x"0FECF",x"0FE8C",x"0FE49",x"0FE27",
									 x"0FE06",x"10001",x"0FDE6",x"0FDC6",x"0FDA5",x"10001",x"0FD85",x"0FD64",x"0FD24",x"0F503",
									 x"0F4E3",x"0F4A3",x"0F483",x"0F442",x"0F403",x"0EC88",x"0F5F2",x"0F719",x"0F77D",x"0F7DF",
									 x"0FFDF",x"0FFFF",x"1000E",x"0FFFF",x"10010",x"0FFDE",x"0FF7B",x"0F6D8",x"0F5B1",x"0EC47",
									 x"0EC23",x"0F441",x"0F483",x"0FCC4",x"0FCE3",x"0F524",x"0FD44",x"0FD64",x"0FD84",x"0FDA5",
									 x"10001",x"0FDC5",x"0FDE6",x"0FE06",x"10001",x"0FE27",x"0FE69",x"0FEAD",x"0FEB0",x"10000",
									 x"0FEAF",x"0FECF",x"100A4",x"0FED0",x"0FECF",x"0FE8C",x"0FE49",x"0FE27",x"0FE06",x"10001",
									 x"0FDE6",x"10000",x"0FDA5",x"10001",x"0F585",x"0FD65",x"0FD44",x"0FD03",x"0F4E3",x"0F4C4",
									 x"0F4A3",x"0F442",x"0F422",x"0EC46",x"0F58E",x"0F6B7",x"0F75C",x"0FFDF",x"10000",x"0FFFF",
									 x"1000E",x"0FFFF",x"1000F",x"0FFDF",x"0FFDE",x"0FF19",x"0EE13",x"0ED2D",x"0EC25",x"0EC43",
									 x"0EC62",x"0F4A3",x"0F4E3",x"0F503",x"0FD24",x"0FD64",x"0FD85",x"10000",x"0FDA5",x"10000",
									 x"0FDC5",x"0FDC6",x"0FDE6",x"0FE06",x"10001",x"0FE48",x"0FE6A",x"0FEAD",x"0FECF",x"10000",
									 x"0FECE",x"0FECF",x"10000",x"0FEEF",x"0FECF",x"100A3",x"0FEAD",x"0FE6A",x"0FE48",x"0FE26",
									 x"0FE06",x"10000",x"0FDE7",x"0FDE6",x"0FDC5",x"0FDA5",x"10000",x"0FD85",x"10000",x"0FD64",
									 x"0FD24",x"0FD04",x"0F4E4",x"0F4A3",x"0F463",x"0F422",x"0EC24",x"0ED0B",x"0EDD2",x"0F6FA",
									 x"0FFDF",x"0FFBE",x"0FFDE",x"0FFFF",x"1000D",x"0FFFF",x"1000F",x"0F7DF",x"0FFBE",x"0F6D8",
									 x"0E56F",x"0ECA9",x"0EC04",x"0F443",x"0F462",x"0FCC3",x"0FD03",x"0F523",x"0F544",x"0FD65",
									 x"0FD85",x"10000",x"0FDA5",x"0FDC5",x"10000",x"0FDC6",x"0FDE6",x"0FE06",x"10000",x"0FE27",
									 x"0FE48",x"0FE8B",x"0FEAD",x"0FECF",x"10000",x"0FECE",x"10000",x"0FECF",x"1002E",x"0FEEF",
									 x"0FECF",x"10071",x"0FECE",x"0FECF",x"10000",x"0FEAE",x"0FE8B",x"0FE49",x"0FE27",x"0FE06",
									 x"10000",x"0FDE7",x"0FDE6",x"10000",x"0FDC5",x"0FDA5",x"10000",x"0FD85",x"0FD64",x"0FD24",
									 x"0FD04",x"0F4E3",x"0F4C3",x"0F483",x"0F442",x"0EC24",x"0EC88",x"0E52E",x"0F698",x"0FF9E",
									 x"0F7BE",x"0FFDF",x"0FFFF",x"1000D",x"0FFFF",x"1000F",x"0F7DF",x"0F79E",x"0F696",x"0ECEB",
									 x"0F466",x"0EC23",x"0F462",x"0F482",x"0FCC4",x"0FD04",x"0FD24",x"0F544",x"0FD65",x"0FD85",
									 x"0FDA5",x"10000",x"0FDC6",x"10000",x"0FDE6",x"0FE06",x"10001",x"0FE27",x"0FE49",x"0FE8B",
									 x"0FEAD",x"0FECF",x"10000",x"0FECE",x"10002",x"0FECF",x"0FECE",x"10029",x"0FECF",x"0FEEF",
									 x"10000",x"0FECE",x"10000",x"0FECF",x"10001",x"0FECE",x"1003A",x"0FECF",x"10003",x"0FECE",
									 x"1002D",x"0FECF",x"0FEAE",x"0FE8C",x"0FE69",x"0FE47",x"0FE26",x"0FE06",x"0FDE7",x"0FDE6",
									 x"10000",x"0FDC6",x"0FDC5",x"0FDA5",x"0FD85",x"0FD65",x"0FD44",x"10000",x"0F503",x"0F4C3",
									 x"0F4A3",x"0F462",x"0EC23",x"0EC66",x"0ECCA",x"0F634",x"0FF7C",x"0F7BE",x"0FFFF",x"1000E",
									 x"0FFFF",x"1000E",x"0F7DE",x"0F7BE",x"0F75B",x"0F613",x"0EC68",x"0F424",x"0F443",x"0F482",
									 x"0F4A3",x"0FCE4",x"0FD04",x"0FD44",x"0FD64",x"0FD85",x"0FDA5",x"10000",x"0FDC5",x"0FDC6",
									 x"10000",x"0FDE6",x"0FE06",x"0FE27",x"0FE26",x"0FE27",x"0FE6A",x"0FEAC",x"0FECE",x"1002F",
									 x"0FEEF",x"0FECE",x"0FEEF",x"10002",x"0FEEE",x"10002",x"0FEEF",x"0FECE",x"10000",x"0FEEF",
									 x"0FECE",x"1002D",x"0FEEF",x"10001",x"0FECE",x"0FEEF",x"10001",x"0FECE",x"0FEEF",x"0FECF",
									 x"10002",x"0FEEF",x"0FECE",x"10000",x"0FEEF",x"0FECE",x"0FEEF",x"10000",x"0FECE",x"10027",
									 x"0FEAF",x"10000",x"0FEAD",x"0FE6A",x"0FE27",x"0FE26",x"0FE06",x"0FDE6",x"10002",x"0FDC6",
									 x"0FDA5",x"10000",x"0FD85",x"0FD64",x"0FD44",x"0F523",x"0F4E3",x"0F4C3",x"0F482",x"0F443",
									 x"0F444",x"0EC67",x"0ED90",x"0FF1A",x"0EF7D",x"0FFFF",x"1000E",x"0FFFF",x"1000E",x"0F7BE",
									 x"0F77D",x"0EEB8",x"0ED6F",x"0EC25",x"0F423",x"0F463",x"0FCA2",x"0F4E3",x"0F504",x"0FD24",
									 x"0FD44",x"0FD64",x"0FD85",x"0FDA5",x"0FDC5",x"0FDC6",x"0FDE6",x"10001",x"0FE06",x"0FE27",
									 x"0FE26",x"0FE47",x"0FE8B",x"0FEAC",x"0FEAD",x"0FECE",x"10000",x"0FEAE",x"0FECE",x"1002A",
									 x"0FEEE",x"10001",x"0FECE",x"10004",x"0FEEE",x"10001",x"0FECE",x"1002C",x"0FEAE",x"0FECE",
									 x"10001",x"0FEEE",x"0FECE",x"10000",x"0FEEE",x"10002",x"0FECE",x"10000",x"0FEAE",x"0FECF",
									 x"10000",x"0FECE",x"0FEEE",x"10000",x"0FECE",x"10029",x"0FEAE",x"0FECD",x"0FECE",x"0FEAF",
									 x"10000",x"0FEAD",x"0FE8B",x"0FE48",x"0FE26",x"0FE06",x"10000",x"0FDE6",x"10001",x"0FDC6",
									 x"10000",x"0FDA5",x"0FD85",x"0FD65",x"0FD64",x"0FD44",x"0F503",x"0F4E3",x"0F4A3",x"0F463",
									 x"0F423",x"0EC24",x"0ED0C",x"0F676",x"0EF5C",x"0F7DF",x"10000",x"0FFFF",x"1000C",x"0FFFF",
									 x"1000D",x"0FFDF",x"0F7BF",x"0F75C",x"0EE55",x"0ED0C",x"0EC24",x"0F423",x"0F463",x"0F4C2",
									 x"0F503",x"0F524",x"0F544",x"0FD64",x"0FD85",x"10000",x"0FDA5",x"0FDC6",x"0FDE6",x"10000",
									 x"0FE06",x"10001",x"0FE27",x"0FE26",x"0FE48",x"0FE6B",x"0FEAD",x"10000",x"0FEAE",x"10003",
									 x"0FECE",x"10026",x"0FEAE",x"0FECE",x"10002",x"0F68C",x"0F68D",x"0EE6C",x"0EE4C",x"10000",
									 x"0F68C",x"0FEAD",x"0FECD",x"0FECE",x"0FEEE",x"0FECE",x"1002C",x"0FEAE",x"0FECE",x"10002",
									 x"0FEEE",x"0FECE",x"10000",x"0FEAE",x"0F6AD",x"0EE6C",x"0EE4C",x"0EE4D",x"0F66D",x"0F68D",
									 x"0FEAE",x"0FECE",x"0FEEE",x"0FECE",x"10029",x"0FEAE",x"0FEAD",x"0FEAE",x"10001",x"0FEAD",
									 x"0FE8B",x"0FE48",x"0FE26",x"10000",x"0FE07",x"0FE06",x"10000",x"0FDE6",x"10000",x"0FDC6",
									 x"0FDA5",x"10000",x"0FD85",x"0FD65",x"0FD44",x"0F524",x"0FCE4",x"0F4A3",x"0F483",x"0F422",
									 x"0F403",x"0ECCA",x"0EE14",x"0F75C",x"0F7DE",x"0F7DF",x"0FFFF",x"1000C",x"0FFFF",x"1000C",
									 x"0FFDF",x"0FFDE",x"0F7BD",x"0F75B",x"0F5F2",x"0F488",x"0F444",x"0EC43",x"0F483",x"0FCC3",
									 x"0FCE4",x"0FD24",x"0FD44",x"0FD64",x"0FD85",x"0FDA5",x"0FDC5",x"0FDE6",x"10002",x"0FE06",
									 x"10000",x"0FE26",x"0FE27",x"0FE48",x"0FE8C",x"0FEAC",x"0FEAD",x"10000",x"0FEAE",x"10000",
									 x"0FEAD",x"0FECE",x"10003",x"0FECD",x"1001E",x"0FECE",x"10001",x"0FECD",x"0FEEE",x"0FEEF",
									 x"0FEEE",x"0F68D",x"0E60C",x"0D54A",x"0C4E9",x"0BCC9",x"0BCC8",x"0C4E9",x"0CD29",x"0DDCC",
									 x"0F68D",x"0F6CD",x"0FEEF",x"10001",x"0FECD",x"10000",x"0FEAD",x"0FECE",x"0FECD",x"10002",
									 x"0FEAD",x"0FECD",x"10003",x"0FECE",x"10004",x"0FECD",x"1000A",x"0FECE",x"10008",x"0FEAE",
									 x"10000",x"0FECE",x"10000",x"0FECD",x"10000",x"0FF0E",x"0FEED",x"10000",x"0F6AD",x"0E62D",
									 x"0CD4A",x"0BCE9",x"0BCC8",x"0BCA8",x"0C4E9",x"0CD4A",x"0E5EB",x"0F6AE",x"0FEEE",x"10001",
									 x"0FECE",x"10001",x"0FECD",x"1000C",x"0FECE",x"10003",x"0FECD",x"1000E",x"0FEAD",x"10001",
									 x"0FECD",x"0FEAD",x"0FEAE",x"10002",x"0FE8B",x"0FE48",x"0FE26",x"0FE06",x"0FE07",x"0FE06",
									 x"10000",x"0FDE6",x"10000",x"0FDC6",x"0FDC5",x"0FDA5",x"0FD85",x"10000",x"0FD64",x"0FD24",
									 x"0FD03",x"0F4C3",x"0F483",x"0F463",x"0EC43",x"0EC67",x"0F5B0",x"0F71A",x"0F79E",x"0FFDE",
									 x"0FFDF",x"10000",x"0FFFF",x"1000A",x"0FFFF",x"1000C",x"0FFDF",x"0FFBE",x"0F77C",x"0F6D8",
									 x"0ED6F",x"0EC26",x"0F423",x"0EC63",x"0F483",x"0FCE4",x"0FD04",x"0FD24",x"0FD44",x"0FD85",
									 x"10000",x"0FDA5",x"0FDC5",x"0FDE6",x"10000",x"0FE06",x"10002",x"0FE26",x"0FE27",x"0FE48",
									 x"0FE8B",x"0FEAC",x"0FEAD",x"10004",x"0FECD",x"10020",x"0FEAD",x"10001",x"0FECD",x"10000",
									 x"0FEED",x"0FECD",x"0EE4C",x"0DDCB",x"0BCE9",x"0A3E7",x"08B25",x"07AA3",x"07282",x"10000",
									 x"072A3",x"082E4",x"09BC7",x"0B4A9",x"0C52A",x"0E60C",x"0F6AE",x"0FEEE",x"0FECD",x"10000",
									 x"0F68D",x"0FECD",x"10003",x"0FEAD",x"10000",x"0FECD",x"10014",x"0FECE",x"10007",x"0FEAE",
									 x"0FEAD",x"10000",x"0FECE",x"0FECD",x"0FEED",x"10000",x"0FECE",x"0E64C",x"0CD4A",x"0BCC9",
									 x"09BC7",x"08304",x"07AA3",x"07281",x"07282",x"07AC3",x"08304",x"09BC6",x"0BCC9",x"0D58B",
									 x"0EE2C",x"0FECD",x"0FEEE",x"0FECD",x"0FEAD",x"0FECD",x"10021",x"0FEAD",x"10004",x"0FEAE",
									 x"10001",x"0FE8C",x"0FE49",x"0FE27",x"0FE07",x"10000",x"0FE06",x"10001",x"0FDE6",x"10000",
									 x"0FDC6",x"0FDA5",x"0FD85",x"10000",x"0FD64",x"0FD44",x"0FD03",x"0F4E4",x"0F4A3",x"0F463",
									 x"0F443",x"0EC46",x"0F52D",x"0F6B8",x"0F75C",x"0FFBE",x"0F7DF",x"0FFDF",x"0FFFE",x"0FFFF",
									 x"10009",x"0FFFF",x"1000B",x"0FFDF",x"10000",x"0FFBE",x"0F71A",x"0EE55",x"0ED0C",x"0EC05",
									 x"0F443",x"0F463",x"0F4A3",x"0FCE4",x"0FD24",x"0FD44",x"0FD64",x"0FD85",x"0FDA5",x"10000",
									 x"0FDC6",x"0FDE6",x"10000",x"0FE06",x"10001",x"0FE26",x"0FE27",x"10000",x"0FE49",x"0FE8C",
									 x"0FEAD",x"1002A",x"0FEAC",x"0FEAD",x"0FECE",x"0EE4C",x"0BCE8",x"093A5",x"06A22",x"05181",
									 x"10000",x"05180",x"10002",x"05140",x"05141",x"059A1",x"07282",x"0AC47",x"0E5EC",x"0F6AD",
									 x"0FEED",x"10000",x"0FECD",x"10000",x"0FEAD",x"10023",x"0FECD",x"0FEAD",x"10001",x"0FECD",
									 x"0FEED",x"0F68C",x"0E5EC",x"0B488",x"07283",x"059C1",x"05161",x"10000",x"05181",x"05160",
									 x"051A0",x"05180",x"05161",x"10000",x"06A02",x"09345",x"0BCA8",x"0E60B",x"0F6AE",x"0FECE",
									 x"0FECD",x"10000",x"0FEAD",x"10029",x"0FE8C",x"0FE49",x"0FE27",x"10000",x"0FE07",x"0FE26",
									 x"0FE06",x"10001",x"0FDE6",x"0FDC6",x"0FDA5",x"10000",x"0FD85",x"0FD64",x"0FD44",x"0FD04",
									 x"0FCE4",x"0F4A3",x"0F463",x"0F443",x"0F425",x"0ECCB",x"0F635",x"0F6FA",x"0F79D",x"0F7DF",
									 x"0FFDF",x"0FFDE",x"0FFFF",x"10009",x"0FFFF",x"1000B",x"0FFDF",x"10000",x"0FFBE",x"0F6D9",
									 x"0F5D1",x"0F4CA",x"0EC04",x"0F443",x"0F483",x"0F4C3",x"0FD04",x"0FD24",x"0FD44",x"0FD84",
									 x"0FDA5",x"10000",x"0FDC5",x"0FDC6",x"0FDE6",x"10000",x"0FE06",x"0FE26",x"10001",x"0FE27",
									 x"10000",x"0FE49",x"0FE6C",x"0FEAD",x"0FECD",x"10000",x"0FEAD",x"10009",x"0FEAC",x"10004",
									 x"0FEAD",x"10011",x"0FEAC",x"0FEAD",x"10001",x"0FEAC",x"0FECD",x"0FEAD",x"0EE4D",x"0C4E9",
									 x"09386",x"07284",x"05981",x"04900",x"04960",x"05180",x"059A0",x"10001",x"05140",x"04940",
									 x"05140",x"05980",x"08304",x"0BCA8",x"0DDCA",x"0F68C",x"0FEED",x"0FECD",x"10000",x"0FEAD",
									 x"0FECD",x"0FEAC",x"10001",x"0FEAD",x"1001F",x"0FECD",x"10001",x"0FEEE",x"0F6AD",x"0DDCB",
									 x"0BCC9",x"08B25",x"061C2",x"05140",x"04900",x"05160",x"05180",x"10001",x"05160",x"05161",
									 x"04920",x"05160",x"07262",x"09344",x"0BCE8",x"0EE2C",x"0FEAD",x"0FEED",x"0FECD",x"0FEAD",
									 x"10004",x"0FEAC",x"0FEAD",x"10007",x"0FEAC",x"10003",x"0FEAD",x"10014",x"0FE8C",x"0FE6A",
									 x"0FE47",x"0FE27",x"10000",x"0FE26",x"0FE06",x"10000",x"0FDE6",x"10000",x"0FDC6",x"0FDC5",
									 x"0FDA5",x"0FD85",x"0FD84",x"0FD44",x"0FD24",x"0FD04",x"0F4C3",x"0F483",x"0F443",x"0F424",
									 x"0EC89",x"0F5D1",x"0F6B8",x"0FF9D",x"0F7DF",x"0FFDF",x"0FFDE",x"0FFFF",x"10009",x"0FFFF",
									 x"1000B",x"0FFDF",x"0F7BE",x"0FFBE",x"0F697",x"0F56E",x"0F487",x"0EC03",x"0F463",x"0F4A2",
									 x"0F4E3",x"0FD04",x"0FD44",x"0FD64",x"0FD84",x"0FDA5",x"10000",x"0FDC6",x"0FDE6",x"10000",
									 x"0FE06",x"10000",x"0FE26",x"10001",x"0FE27",x"0FE48",x"0FE69",x"0FE8C",x"0FEAD",x"0FECD",
									 x"0FEAD",x"0FEAC",x"10024",x"0FE8C",x"0FEAC",x"10000",x"0FECD",x"0EE2C",x"0C50A",x"08B05",
									 x"061A1",x"05981",x"059C1",x"061E1",x"06200",x"06A20",x"06A00",x"10000",x"06A01",x"10000",
									 x"061E1",x"059C1",x"05980",x"059A0",x"07AA3",x"0A3C5",x"0DDAB",x"0FEAD",x"0FEEE",x"0FECD",
									 x"0FEAD",x"0FECD",x"0FEAC",x"0FEAD",x"0FEAC",x"10017",x"0FEAD",x"10005",x"0FEAC",x"10001",
									 x"0FEED",x"10000",x"0FECD",x"0DDCB",x"0AC27",x"07AC3",x"059A0",x"10001",x"061C1",x"06201",
									 x"06A01",x"06A00",x"10000",x"06A01",x"06201",x"061C0",x"059C0",x"059A0",x"10000",x"082C3",
									 x"0BCC9",x"0E60B",x"0FECD",x"10000",x"0FECC",x"10000",x"0FEAC",x"0FECC",x"0FEAC",x"10022",
									 x"0FEAD",x"10001",x"0FE8C",x"0FE6A",x"0FE48",x"0FE27",x"10000",x"0FE26",x"0FE06",x"10001",
									 x"0FDE6",x"10000",x"0FDC5",x"0FDA5",x"10000",x"0FD84",x"0FD44",x"0FD24",x"0FD04",x"0F4E3",
									 x"0F4A3",x"0F463",x"0F423",x"0EC67",x"0F54D",x"0F675",x"0FF7C",x"0FFDF",x"10000",x"0FFDE",
									 x"0FFFF",x"10009",x"0FFFF",x"1000B",x"0FFDF",x"0F7BE",x"0F79D",x"0EE55",x"0ED0B",x"0F446",
									 x"0EC03",x"0F482",x"0F4C2",x"0F4E3",x"0FD24",x"0FD44",x"0FD64",x"0FDA4",x"0FDA5",x"10000",
									 x"0FDC6",x"0FDE6",x"0FE06",x"10000",x"0FE26",x"10002",x"0FE47",x"0FE48",x"0FE6A",x"0FE8C",
									 x"0FEAD",x"0FEAC",x"10025",x"0FECC",x"0FEAD",x"0FECD",x"0FECC",x"0F66B",x"0C4E8",x"08B24",
									 x"061C1",x"05180",x"061C0",x"06A00",x"07241",x"07242",x"07241",x"07261",x"10000",x"07241",
									 x"10000",x"07221",x"06A21",x"06201",x"059A1",x"10000",x"07241",x"0AC06",x"0DDCA",x"0FECD",
									 x"10000",x"0FEAC",x"0FEAD",x"0FEAC",x"0FECC",x"0FEAC",x"1001C",x"0FE8C",x"0FEAC",x"10001",
									 x"0FECC",x"0FEED",x"0FECC",x"0E5EA",x"0AC26",x"07261",x"059A0",x"10000",x"061E1",x"06A01",
									 x"07241",x"10000",x"07261",x"10000",x"07241",x"07A42",x"07241",x"10000",x"06A21",x"059C1",
									 x"05981",x"061C0",x"08B03",x"0BCC7",x"0EE4B",x"0FECD",x"0FECC",x"0FECD",x"0FEAC",x"10026",
									 x"0FEAD",x"0FE8C",x"0FE6A",x"0FE48",x"10000",x"0FE27",x"0FE26",x"10000",x"0FE06",x"10001",
									 x"0FDE6",x"0FDC6",x"0FDA5",x"10000",x"0FD85",x"0FD64",x"0FD44",x"0FD24",x"0F504",x"0F4C3",
									 x"0F483",x"0F443",x"0EC45",x"0E4EA",x"0EE13",x"0F75C",x"0FFBE",x"0F7BF",x"0FFDF",x"0FFFF",
									 x"10009",x"0FFFF",x"1000B",x"0F7BF",x"0F7BD",x"0FF5B",x"0EE12",x"0ECA9",x"0F424",x"0F443",
									 x"0F483",x"0F4A3",x"0FD03",x"0FD24",x"0FD44",x"0FD64",x"0FDA5",x"10001",x"0FDC6",x"0FDE6",
									 x"0FE06",x"10000",x"0FE26",x"10002",x"0FE47",x"0FE48",x"0FE6A",x"0FE8C",x"0FEAC",x"10026",
									 x"0FECB",x"0FEAC",x"0FEAD",x"0FEAC",x"0DDCA",x"0AC26",x"06A21",x"05980",x"061E0",x"06A20",
									 x"07240",x"07A41",x"07A61",x"10005",x"07241",x"07201",x"069E0",x"05980",x"061C0",x"08304",
									 x"0C4E8",x"0F6AD",x"0FECD",x"0FEEC",x"0FEAC",x"0FECC",x"0FEAC",x"1001F",x"0FEAD",x"0FEAC",
									 x"0FECC",x"0FEED",x"0F68C",x"0CD49",x"09345",x"061C1",x"05980",x"06A01",x"07221",x"07241",
									 x"07A61",x"10005",x"07A41",x"07221",x"06A00",x"069E1",x"05980",x"06A00",x"09BC5",x"0DDAA",
									 x"0F6AD",x"0FECD",x"0FEAC",x"10000",x"0FEAB",x"0FEAC",x"10025",x"0FE8D",x"0FE6A",x"0FE48",
									 x"0FE27",x"10001",x"0FE26",x"10000",x"0FE06",x"10000",x"0FDE6",x"0FDC6",x"0FDC5",x"10000",
									 x"0FDA5",x"0FD85",x"0FD64",x"0FD44",x"0FD04",x"0F4C3",x"0F4A2",x"0F462",x"0EC45",x"0ECA9",
									 x"0F5D1",x"0FF3A",x"0F7BD",x"0F7DE",x"0FFDF",x"0FFFF",x"10009",x"0FFFF",x"1000A",x"0F7FF",
									 x"0F7BE",x"0F77C",x"0F6F8",x"0EDB0",x"0EC88",x"0F423",x"0F463",x"0F4A3",x"0F4C3",x"0FD04",
									 x"0FD24",x"0FD44",x"0FD64",x"0FDA5",x"10001",x"0FDC6",x"0FDE6",x"0FE06",x"10000",x"0FE26",
									 x"10001",x"0FE46",x"0FE47",x"0FE48",x"0FE6A",x"0FE8C",x"0FEAC",x"10000",x"0FEAB",x"0FEAC",
									 x"10023",x"0FECB",x"0FECC",x"0FECD",x"0EE4C",x"0B487",x"08B03",x"061E0",x"061A0",x"07201",
									 x"07241",x"07A61",x"07A81",x"082A1",x"08281",x"10002",x"082A2",x"07A81",x"07A61",x"10000",
									 x"07220",x"061A0",x"10000",x"07241",x"09BC5",x"0DDCA",x"0F68C",x"0FEED",x"0FEAB",x"0FEAC",
									 x"10020",x"0FEAD",x"0FEAC",x"0FEEC",x"0F6AC",x"0DDCA",x"0AC06",x"07262",x"061A1",x"061A0",
									 x"07221",x"07A41",x"07A61",x"07A81",x"08281",x"10000",x"082A1",x"10001",x"08281",x"10000",
									 x"07A61",x"07220",x"07221",x"061C0",x"10000",x"07AC2",x"0AC66",x"0EE4C",x"0FECD",x"0FEAD",
									 x"0FEAC",x"0FEAB",x"0FEAC",x"10025",x"0FE8C",x"0FE6A",x"0FE48",x"0FE47",x"0FE27",x"10001",
									 x"0FE26",x"0FE06",x"10000",x"0FDE6",x"0FDC6",x"0FDC5",x"10000",x"0FDA5",x"0FD85",x"0FD64",
									 x"0FD44",x"0FD04",x"0F4E3",x"0F4C2",x"0F483",x"0EC44",x"0EC67",x"0ED6F",x"0F6D8",x"0F77C",
									 x"0F7BE",x"0F7DF",x"0FFFF",x"10009",x"0FFFF",x"1000A",x"0F7DF",x"0F7BE",x"0F75B",x"0F696",
									 x"0ED2D",x"0EC66",x"0F422",x"0F483",x"0F4C3",x"0FD04",x"10000",x"0FD24",x"0FD64",x"0FD84",
									 x"0FDA5",x"0FDC5",x"0FDC6",x"10000",x"0FDE6",x"0FE06",x"10000",x"0FE26",x"10001",x"0FE46",
									 x"0FE47",x"0FE48",x"0FE6A",x"0FE8C",x"0FEAC",x"10000",x"0FE8B",x"0FE8C",x"0FEAC",x"10018",
									 x"0FE8C",x"10003",x"0FEAC",x"10001",x"0FE8C",x"0FEAC",x"0FEAB",x"0FECB",x"0FEAC",x"0DDCB",
									 x"08B23",x"061E0",x"10000",x"06A00",x"07A62",x"07A81",x"08281",x"082A1",x"10000",x"08AA1",
									 x"10001",x"08AC1",x"10000",x"082A1",x"082A2",x"08282",x"07A61",x"07221",x"069E1",x"059A0",
									 x"07AA2",x"0BCC7",x"0E5EA",x"0FEED",x"0FECC",x"0FEAC",x"10003",x"0FE8C",x"10007",x"0FEAC",
									 x"10004",x"0FE8C",x"1000A",x"0FEAC",x"10002",x"0FEED",x"0E62B",x"0BCC8",x"082E3",x"059A0",
									 x"061C1",x"07201",x"07A61",x"08281",x"10000",x"082A1",x"08AC1",x"10002",x"08AA1",x"082A1",
									 x"10000",x"08281",x"07A61",x"10000",x"07201",x"061C1",x"061E1",x"082E2",x"0D58A",x"0FEAC",
									 x"10001",x"0FEAB",x"0FEAC",x"10022",x"0FE8C",x"0FEAC",x"10000",x"0FE8C",x"0FE6A",x"0FE48",
									 x"0FE27",x"10004",x"0FE06",x"0FDE6",x"0FDC6",x"0FDC5",x"10000",x"0FDA5",x"0FD85",x"0FD65",
									 x"0FD44",x"0F504",x"0F4E4",x"0F4E3",x"0F482",x"0F423",x"0EC25",x"0ED0C",x"0F655",x"0F73B",
									 x"0F7BE",x"0F7DF",x"0FFFF",x"10009",x"0FFFF",x"10009",x"0FFDF",x"0F7DF",x"0F7BE",x"0F73A",
									 x"0F633",x"0ECEB",x"0EC45",x"0F442",x"0F482",x"0F4C3",x"0F504",x"0FD04",x"0FD44",x"0FD65",
									 x"0FD85",x"0FDA5",x"0FDC5",x"0FDC6",x"0FDE6",x"0FE06",x"10001",x"0FE26",x"10001",x"0FE47",
									 x"10000",x"0FE48",x"0FE6A",x"0FE8B",x"0FEAC",x"10000",x"0FE8B",x"0FEAC",x"10019",x"0FE8C",
									 x"10006",x"0FEAC",x"10000",x"0FEAB",x"10000",x"0EE4B",x"0CD0A",x"07242",x"05980",x"06A01",
									 x"07A41",x"08282",x"08281",x"082A1",x"08AC1",x"08AE2",x"092E1",x"10002",x"08AE1",x"08AC1",
									 x"10000",x"082A1",x"10000",x"07A61",x"07221",x"05980",x"06A21",x"0A3E5",x"0CD49",x"0FEAC",
									 x"0FECC",x"0FEAC",x"10021",x"0FECC",x"0FECD",x"0D589",x"0A3E6",x"07241",x"05980",x"07201",
									 x"07A41",x"08281",x"10000",x"082A1",x"08AC1",x"10000",x"092E1",x"10001",x"08AE1",x"08AC1",
									 x"08AC2",x"082A1",x"08281",x"07A61",x"10000",x"07223",x"061A1",x"06A21",x"0BCC8",x"0EE4B",
									 x"0F68C",x"0FEAC",x"0FE8B",x"0FEAC",x"10001",x"0FE8C",x"10003",x"0FEAC",x"1001A",x"0FE8C",
									 x"0FEAC",x"10000",x"0FE8C",x"0FE6A",x"0FE68",x"0FE48",x"0FE28",x"0FE27",x"10001",x"0FE26",
									 x"0FE06",x"10000",x"0FDE6",x"0FDE5",x"10000",x"0FDC5",x"0FD85",x"0FD65",x"0FD45",x"0FD25",
									 x"0F504",x"0F503",x"0F482",x"0F443",x"0F424",x"0ECC9",x"0F5F2",x"0F71A",x"0F7BE",x"0F7DF",
									 x"0FFFF",x"0FFDF",x"0FFFF",x"10007",x"0FFFF",x"10009",x"0FFDF",x"0F7DF",x"0F7BE",x"0F71A",
									 x"0EDD1",x"0ECA9",x"0EC44",x"0FC42",x"0F4A3",x"0F4C4",x"0F504",x"0FD24",x"0FD44",x"0FD65",
									 x"0FD85",x"0FDA5",x"0FDC5",x"0FDE6",x"10000",x"0FE06",x"10001",x"0FE26",x"10001",x"0FE47",
									 x"10000",x"0FE48",x"0FE69",x"0FE8B",x"10000",x"0FE8C",x"10000",x"0FE8B",x"0FEAB",x"0FEAC",
									 x"10017",x"0FE8C",x"10007",x"0FEAC",x"0FEAB",x"0F68B",x"0DDAA",x"0B468",x"07221",x"061C0",
									 x"07221",x"07A81",x"08281",x"082A1",x"08AC1",x"08AE1",x"09301",x"09302",x"09B02",x"09302",
									 x"10000",x"092E2",x"10000",x"092C2",x"08AA2",x"082A1",x"08281",x"07A42",x"061C1",x"07221",
									 x"09365",x"0BCC8",x"0F66C",x"0FECB",x"0FEAC",x"10000",x"0FE8B",x"10000",x"0FE8C",x"10002",
									 x"0FEAC",x"10004",x"0FEAB",x"10004",x"0FEAC",x"10004",x"0FE8C",x"10004",x"0FEAB",x"0FEAC",
									 x"10000",x"0FECC",x"0F68C",x"0C508",x"09365",x"07241",x"061A0",x"07A41",x"08261",x"08AA1",
									 x"10000",x"08AC1",x"092C1",x"092E1",x"10003",x"092E2",x"10000",x"08AC1",x"08AA1",x"08281",
									 x"07A61",x"07222",x"061E1",x"06A21",x"0AC26",x"0DDAA",x"0F66B",x"0FECC",x"0FEAB",x"10000",
									 x"0FE8C",x"0FEAC",x"0FE8C",x"10004",x"0FEAC",x"10018",x"0FE8C",x"10001",x"0FEAC",x"0FE8B",
									 x"0FE89",x"0FE48",x"10000",x"0FE28",x"0FE47",x"0FE27",x"10000",x"0FE26",x"0FE06",x"10000",
									 x"0FDE6",x"10000",x"0FDE5",x"0FDA5",x"0FD85",x"0FD65",x"10000",x"0FD25",x"0F504",x"0F503",
									 x"0F4A3",x"0F443",x"0F423",x"0EC87",x"0ED6F",x"0F6F9",x"0F79E",x"0F7DF",x"0FFFF",x"0FFDF",
									 x"0FFFF",x"10007",x"0FFFF",x"10009",x"0FFDF",x"0F7BF",x"0F77D",x"0F6D8",x"0E56F",x"0E487",
									 x"0F423",x"0F442",x"0FCA3",x"0FCC4",x"0FD04",x"0FD44",x"0FD65",x"0FD85",x"0FDA5",x"0FDC5",
									 x"10000",x"0FDE6",x"0FE06",x"10002",x"0FE26",x"10001",x"0FE47",x"10000",x"0FE48",x"0FE69",
									 x"0FE8B",x"10000",x"0FE8C",x"10000",x"0FEAB",x"10000",x"0FEAC",x"0FE8C",x"0FEAC",x"0FE8C",
									 x"1001D",x"0FEAC",x"0FEAB",x"0F66C",x"0CD29",x"09BC5",x"06A20",x"06A00",x"07A41",x"08282",
									 x"08AA1",x"08AC1",x"10000",x"092E1",x"09301",x"09B02",x"10002",x"09302",x"10000",x"092E3",
									 x"08AC2",x"08AC1",x"082A1",x"07A62",x"07201",x"10000",x"082E3",x"0AC26",x"0EE2A",x"0FECB",
									 x"0FECC",x"0FEAC",x"0FE8B",x"1000B",x"0FE8A",x"10002",x"0FE8B",x"1000C",x"0FEAC",x"0FECD",
									 x"0FECC",x"0EE4B",x"0B486",x"08303",x"06A21",x"06A00",x"07A61",x"08281",x"08AC1",x"092C1",
									 x"092E2",x"09B02",x"10001",x"09B01",x"10001",x"09302",x"092E2",x"08AC1",x"10000",x"08AA1",
									 x"08281",x"07A42",x"06A01",x"06A20",x"09384",x"0C508",x"0EE4B",x"0FECC",x"0FEAB",x"0FE8B",
									 x"0FE8C",x"10011",x"0FEAC",x"10002",x"0FE8C",x"10004",x"0FEAC",x"10001",x"0FE8C",x"10001",
									 x"0FE8B",x"0FE8C",x"10000",x"0FE8B",x"0FE69",x"0FE48",x"0FE28",x"10000",x"0FE47",x"0FE27",
									 x"10000",x"0FE26",x"0FE06",x"10000",x"0FDE6",x"0FDE5",x"10000",x"0FDC5",x"0FDA5",x"0FD85",
									 x"0FD65",x"0FD24",x"0FD04",x"0F503",x"0F4C3",x"0F463",x"0F423",x"0EC66",x"0ED2D",x"0F6B8",
									 x"0EF7D",x"0F7BF",x"0F7DF",x"0FFFF",x"10008",x"0FFFF",x"10009",x"0FFBE",x"0F79E",x"0F75C",
									 x"0F676",x"0ED0D",x"0EC46",x"0EC44",x"0F462",x"0F4A2",x"0F4E4",x"0F504",x"0FD44",x"0FD65",
									 x"0FD85",x"0FDA5",x"10000",x"0FDC6",x"0FDE6",x"0FE06",x"10001",x"0FE26",x"0FE27",x"0FE26",
									 x"10000",x"0FE46",x"0FE47",x"0FE68",x"0FE89",x"0FE8A",x"0FE8B",x"10002",x"0FEAB",x"0FE8B",
									 x"10010",x"0FEAB",x"10008",x"0FE8B",x"10000",x"0FEAB",x"10001",x"0FE8B",x"0FEAB",x"0FECB",
									 x"0EE6B",x"0BCE7",x"08B03",x"06A21",x"07221",x"07A61",x"082A1",x"08AC1",x"10000",x"092E1",
									 x"09301",x"09B21",x"09B22",x"0A322",x"10000",x"09B22",x"10000",x"09B02",x"092E2",x"10000",
									 x"08AC1",x"08AA1",x"08281",x"07241",x"07201",x"07A82",x"09BA4",x"0DDC9",x"0FEAA",x"0FECB",
									 x"0FE8B",x"0FE6A",x"0FE8A",x"10000",x"0FE6A",x"0FE69",x"10005",x"0FE89",x"1000C",x"0FE69",
									 x"10003",x"0FE6A",x"0FE8A",x"0FECB",x"10000",x"0E5EA",x"0A405",x"07A82",x"06A21",x"07240",
									 x"08281",x"082A1",x"08AC1",x"092E2",x"09AE2",x"09B02",x"09B22",x"0A322",x"10000",x"09B21",
									 x"09B22",x"10000",x"09B02",x"092E1",x"092C1",x"08AC1",x"08AA2",x"08261",x"07241",x"07220",
									 x"082E3",x"0BCA7",x"0EE4B",x"0FECB",x"0FEAB",x"10000",x"0FE8B",x"10015",x"0FEAB",x"10004",
									 x"0FE8B",x"10007",x"0FE8A",x"0FE69",x"0FE68",x"0FE48",x"0FE47",x"10001",x"0FE27",x"10000",
									 x"0FE26",x"0FE06",x"10001",x"0FDE5",x"0FDC5",x"0FDA5",x"0FD84",x"0FD64",x"0FD44",x"0FD23",
									 x"0F503",x"0F4C3",x"0F463",x"0F443",x"0EC45",x"0E4EA",x"0F676",x"0F75C",x"0F79D",x"0FFDF",
									 x"10000",x"0FFFF",x"10007",x"0FFFF",x"10008",x"0FFDF",x"0F7BF",x"0F77D",x"0F71B",x"0F655",
									 x"0ECCB",x"0EC25",x"0F444",x"0F482",x"0F4C2",x"0FD04",x"0F524",x"0FD44",x"0FD65",x"0FD85",
									 x"0FDA5",x"0FDC6",x"10000",x"0FDE6",x"0FE06",x"10001",x"0FE26",x"0FE27",x"0FE26",x"10000",
									 x"0FE46",x"0FE47",x"0FE68",x"0FE89",x"0FE8A",x"0FE8B",x"10001",x"0FEAB",x"0FE8B",x"10021",
									 x"0FEAB",x"0FECC",x"0EE6B",x"0B486",x"07AA2",x"07201",x"07A41",x"08281",x"08AA1",x"092E1",
									 x"10000",x"09301",x"09B02",x"0A322",x"10003",x"09B22",x"10000",x"09B02",x"10000",x"092E1",
									 x"08AC1",x"082A1",x"07A61",x"06A00",x"07221",x"09343",x"0D588",x"0F689",x"0FECA",x"0FE6A",
									 x"0FE49",x"0FE69",x"10000",x"0FE68",x"10002",x"0FE48",x"10000",x"0FE68",x"10014",x"0FE69",
									 x"0FEAA",x"0FEA9",x"0DDA8",x"09BA4",x"07241",x"06A21",x"07A81",x"082A1",x"08AC1",x"092E2",
									 x"10000",x"09B02",x"10000",x"09B22",x"0A322",x"0A342",x"10001",x"0A322",x"09B22",x"09B02",
									 x"092E1",x"092C1",x"08AC1",x"08281",x"07A61",x"07220",x"07A82",x"0B446",x"0EE2B",x"0FECB",
									 x"0FEAB",x"10000",x"0FE8B",x"10024",x"0FE8A",x"0FE69",x"0FE68",x"0FE47",x"10002",x"0FE27",
									 x"10000",x"0FE26",x"0FE06",x"10001",x"0FDE6",x"0FDC5",x"10000",x"0FD85",x"0FD84",x"0FD64",
									 x"0FD24",x"0F503",x"0F4C3",x"0F483",x"0F463",x"0EC44",x"0E4A9",x"0F634",x"0EF1A",x"0EF7D",
									 x"0FFDE",x"0FFDF",x"0FFFF",x"10007",x"0FFFF",x"10008",x"0FFDF",x"0FFBE",x"0EF5D",x"0EED9",
									 x"0F5F2",x"0ECA9",x"0EC24",x"0F463",x"0FCA2",x"0FCE3",x"0FD23",x"0FD44",x"0FD64",x"0FD85",
									 x"10000",x"0FDA5",x"0FDC6",x"0FDE6",x"10000",x"0FE06",x"10001",x"0FE26",x"0FE27",x"10000",
									 x"0FE26",x"0FE46",x"0FE47",x"0FE68",x"0FE89",x"0FE8A",x"10000",x"0FE8B",x"10002",x"0FE8A",
									 x"0FE8B",x"1001F",x"0FEAB",x"0FECC",x"0EE6B",x"0B466",x"07241",x"07221",x"07A61",x"082A1",
									 x"08AC1",x"092E1",x"10000",x"09B01",x"09B22",x"0A322",x"10000",x"0A342",x"10002",x"09B22",
									 x"10000",x"09B02",x"092E1",x"08AE1",x"082A1",x"08281",x"07220",x"06A00",x"08B02",x"0D567",
									 x"0F688",x"0FEC9",x"0FE68",x"0FE47",x"1001C",x"0FE67",x"10000",x"0FEA8",x"0FEA9",x"0D587",
									 x"09363",x"061E0",x"06A00",x"082A2",x"082A1",x"08AE1",x"09302",x"09B02",x"10000",x"09B22",
									 x"0A322",x"0A342",x"10004",x"09B02",x"092E1",x"10000",x"08AC1",x"082A1",x"08281",x"07220",
									 x"07241",x"0AC06",x"0EE2B",x"0FECB",x"0FEAB",x"0FE8B",x"10007",x"0FE8A",x"0FE8B",x"10001",
									 x"0FE8A",x"0FE8B",x"10001",x"0FE8A",x"0FE8B",x"10010",x"0FE8A",x"10002",x"0FE69",x"0FE48",
									 x"0FE47",x"10000",x"0FE27",x"0FE47",x"0FE27",x"10000",x"0FE26",x"0FE06",x"10001",x"0FDE6",
									 x"10000",x"0FDC5",x"0FDA5",x"0FD85",x"0FD64",x"0FD44",x"0F524",x"0F4E4",x"0F483",x"0FC63",
									 x"0F444",x"0E488",x"0EDF2",x"0EEB8",x"0EF5C",x"0F7BE",x"0FFDF",x"0FFFF",x"10007",x"0FFFF",
									 x"10008",x"0FFDF",x"0F7BE",x"0EF5C",x"0EE97",x"0ED90",x"0EC67",x"0EC23",x"0F463",x"0F4A2",
									 x"0FD03",x"0FD24",x"0FD44",x"0FD64",x"0FD85",x"0FDA5",x"10000",x"0FDC6",x"0FDE6",x"0FE06",
									 x"10001",x"0FE27",x"10002",x"0FE47",x"10001",x"0FE67",x"0FE68",x"0FE89",x"0FE6A",x"0FE8A",
									 x"0FE6B",x"0FE6A",x"0FE8A",x"10005",x"0FE8B",x"10004",x"0FE8A",x"10005",x"0FE8B",x"10003",
									 x"0FE8A",x"10005",x"0FE8B",x"10000",x"0FE8A",x"0FE8B",x"0FECB",x"0F66B",x"0AC25",x"06A20",
									 x"07221",x"08281",x"08AA1",x"08AE1",x"092E1",x"09B01",x"09B02",x"0A322",x"10000",x"0A342",
									 x"10004",x"09B22",x"09B02",x"092E1",x"10000",x"08AC1",x"082A2",x"07221",x"061C0",x"08B02",
									 x"0D546",x"0FE88",x"0FEC8",x"0FE67",x"0FE46",x"10000",x"0FE47",x"0FE46",x"0FE47",x"10018",
									 x"0FE46",x"0FE66",x"0FEC8",x"0FEA8",x"0D587",x"09322",x"061C0",x"06A00",x"082A2",x"08AC1",
									 x"092E2",x"10000",x"09B02",x"10000",x"0A322",x"0A342",x"10000",x"0AB42",x"10000",x"0A342",
									 x"10000",x"0A322",x"09B02",x"10000",x"09301",x"092C1",x"08AA1",x"08281",x"07241",x"06A00",
									 x"0A3C5",x"0EE2A",x"0FECB",x"0FEAA",x"0FE8B",x"10000",x"0FE8A",x"10023",x"0FE89",x"0FE68",
									 x"0FE67",x"0FE47",x"10000",x"0FE27",x"0FE47",x"10000",x"0FE27",x"0FE26",x"0FE06",x"10001",
									 x"0FDE6",x"0FDC6",x"0FDC5",x"0FDA5",x"0FD85",x"0FD64",x"0FD44",x"0F524",x"0F504",x"0F4A3",
									 x"0F463",x"0F443",x"0E466",x"0ED90",x"0E656",x"0EF5B",x"0F7BE",x"0F7DF",x"0FFDF",x"0FFFF",
									 x"10006",x"0FFFF",x"10008",x"0FFDE",x"0F7BE",x"0EF3C",x"0EE56",x"0ED4E",x"0EC66",x"0EC23",
									 x"0F463",x"0F4A3",x"0FD04",x"0FD24",x"0FD44",x"0FD64",x"0FD85",x"0FDA5",x"0FDC5",x"0FDC6",
									 x"0FDE6",x"0FE06",x"10000",x"0FE26",x"0FE27",x"10002",x"0FE47",x"10002",x"0FE68",x"10000",
									 x"0FE89",x"0FE8A",x"0FE6A",x"10000",x"0FE8A",x"10020",x"0FE6A",x"0FE8A",x"0FECA",x"0EE6A",
									 x"0A404",x"06A00",x"07221",x"08281",x"08AA1",x"092E1",x"09301",x"09B02",x"09B22",x"0A322",
									 x"0A342",x"0AB42",x"10002",x"0A342",x"10000",x"0A322",x"09B02",x"09B01",x"092E1",x"08AC1",
									 x"082A2",x"07221",x"061A0",x"08AE2",x"0D546",x"0FE88",x"0FEC8",x"0FE67",x"0FE46",x"0FE47",
									 x"10009",x"0FE67",x"10004",x"0FE47",x"1000A",x"0FE46",x"0FE66",x"0FEC8",x"0F6C8",x"0D587",
									 x"09342",x"069E0",x"07220",x"08AC2",x"08AC1",x"092E1",x"09B02",x"09B22",x"09B02",x"0A322",
									 x"0A342",x"10000",x"0AB42",x"0AB62",x"0A342",x"10000",x"0A322",x"09B02",x"10000",x"09B01",
									 x"092E1",x"08AA1",x"08281",x"07A41",x"069E0",x"09BA4",x"0EE2A",x"0FECA",x"0FE89",x"0FE8A",
									 x"10000",x"0FE89",x"0FE8A",x"10022",x"0FE89",x"0FE68",x"0FE67",x"0FE47",x"10003",x"0FE27",
									 x"0FE26",x"0FE06",x"10001",x"0FDE6",x"10000",x"0FDC5",x"0FDA5",x"0FD85",x"0FD65",x"0FD44",
									 x"0F524",x"0F504",x"0F4C3",x"0F483",x"0F442",x"0EC45",x"0ED4E",x"0EE35",x"0F75B",x"0F7DE",
									 x"0F7DF",x"0FFDF",x"0FFFF",x"10006",x"0FFFF",x"10007",x"0FFDF",x"0FFDE",x"0F7BE",x"0EF5C",
									 x"0E635",x"0ED0D",x"0F466",x"0F422",x"0F483",x"0F4C4",x"0FD04",x"0FD25",x"0FD45",x"0FD65",
									 x"0FD85",x"0FDA5",x"0FDC6",x"0FDE6",x"10000",x"0FE06",x"10000",x"0FE26",x"0FE27",x"10000",
									 x"0FE47",x"10004",x"0FE68",x"10000",x"0FE89",x"0FE6A",x"0FE8A",x"0FE6A",x"0FE8A",x"10012",
									 x"0FE6A",x"0FE8A",x"10000",x"0FE6A",x"10000",x"0FE8A",x"10003",x"0FE69",x"10003",x"0FE89",
									 x"0FEA9",x"0EE6A",x"0A404",x"06A00",x"07221",x"08282",x"08AA2",x"092E2",x"09B01",x"09B02",
									 x"0A322",x"10001",x"0AB42",x"10003",x"0A342",x"0A322",x"09B02",x"10000",x"09301",x"08AC2",
									 x"08AA2",x"07221",x"069C0",x"08B02",x"0D546",x"0FE88",x"0FEC8",x"0FE88",x"0FE67",x"10001",
									 x"0FE47",x"10007",x"0FE67",x"10005",x"0FE47",x"1000B",x"0FEC8",x"0F6C8",x"0D587",x"09342",
									 x"069E0",x"07220",x"08AC2",x"08AC1",x"092E1",x"09302",x"09B22",x"0A322",x"10000",x"0AB42",
									 x"10000",x"0AB62",x"10000",x"0A342",x"10000",x"0A322",x"10000",x"09B02",x"10000",x"092E2",
									 x"08AA2",x"08281",x"07A61",x"06A00",x"0A3A3",x"0EE09",x"0FEA9",x"0FE89",x"0FE69",x"10004",
									 x"0FE6A",x"10000",x"0FE8A",x"1001D",x"0FE88",x"0FE67",x"10000",x"0FE47",x"10000",x"0FE27",
									 x"0FE47",x"10000",x"0FE27",x"10000",x"0FE26",x"0FE06",x"10000",x"0FDE6",x"10000",x"0FDC6",
									 x"0FDA6",x"0FD85",x"0FD65",x"0FD45",x"0F524",x"0F504",x"0F4C3",x"0F483",x"0F442",x"0EC44",
									 x"0ED0C",x"0EDF3",x"0F73A",x"0F7DE",x"0F7DF",x"0FFDF",x"0FFFF",x"10006",x"0FFFF",x"10007",
									 x"0FFDF",x"0F7BE",x"10000",x"0F71A",x"0EDF2",x"0ECEA",x"0EC45",x"0F443",x"0F483",x"0FCC4",
									 x"0FD04",x"0FD45",x"0FD65",x"0FD85",x"0FDA5",x"0FDC5",x"0FDC6",x"0FDE6",x"10000",x"0FE06",
									 x"10000",x"0FE26",x"0FE27",x"10000",x"0FE47",x"10005",x"0FE68",x"0FE69",x"10000",x"0FE6A",
									 x"10000",x"0FE8A",x"1000C",x"0FE89",x"10000",x"0FE8A",x"10007",x"0FE89",x"0FE69",x"10002",
									 x"0FE49",x"0FE68",x"10003",x"0FEA8",x"0EE68",x"0AC44",x"07261",x"07241",x"08281",x"08AA2",
									 x"092C2",x"09AE2",x"09B02",x"0A322",x"10000",x"0A342",x"0AB42",x"10003",x"0A342",x"0A322",
									 x"09B22",x"09B02",x"09AE2",x"08AC1",x"082A1",x"07A40",x"07220",x"09322",x"0D587",x"0F6A7",
									 x"0FEE8",x"0FE88",x"0FE47",x"0FE67",x"10000",x"0FE47",x"1001A",x"0FE67",x"0FEC8",x"10000",
									 x"0DDA7",x"09B82",x"07200",x"07241",x"08AC1",x"092C1",x"092C2",x"09B02",x"0A322",x"10000",
									 x"0A342",x"0AB42",x"10000",x"0AB62",x"10000",x"0A342",x"10001",x"0A322",x"09B02",x"09AE2",
									 x"092E2",x"08AC2",x"08281",x"07A41",x"07240",x"0AC04",x"0EE08",x"0FEA9",x"0FE67",x"0FE68",
									 x"10004",x"0FE69",x"10004",x"0FE8A",x"10005",x"0FE89",x"10000",x"0FE8A",x"10000",x"0FE89",
									 x"10009",x"0FE8A",x"10001",x"0FE89",x"0FE68",x"10000",x"0FE67",x"0FE47",x"10003",x"0FE27",
									 x"10001",x"0FE06",x"10001",x"0FDE6",x"10000",x"0FDC6",x"0FDA5",x"10000",x"0FD65",x"0FD44",
									 x"0FD24",x"10000",x"0F4C3",x"0F483",x"0F442",x"0F424",x"0ECEA",x"0EDD1",x"0F6F8",x"0F7BD",
									 x"0F7BE",x"0FFDF",x"0FFFF",x"10006",x"0FFFF",x"10007",x"0FFDF",x"0F7BE",x"0F77D",x"0F6D9",
									 x"0EDB0",x"0ECC9",x"0EC44",x"0F442",x"0F483",x"0FCC4",x"0FD04",x"0FD45",x"0FD65",x"0FD85",
									 x"0FDA5",x"0FDC5",x"0FDC6",x"0FDE6",x"0FE06",x"10001",x"0FE26",x"0FE27",x"10000",x"0FE47",
									 x"10005",x"0FE67",x"0FE68",x"0FE69",x"0FE6A",x"0FE69",x"0FE89",x"0FE8A",x"1000A",x"0FE89",
									 x"10005",x"0FE69",x"10001",x"0FE89",x"10000",x"0FE69",x"0FE68",x"10002",x"0FE48",x"0FE67",
									 x"10000",x"0FE47",x"10000",x"0FE67",x"0FEA8",x"0F688",x"0BCC5",x"08B02",x"07A61",x"08281",
									 x"08AA1",x"092C2",x"09AE2",x"09B02",x"0A322",x"10000",x"0A342",x"0AB42",x"10000",x"0AB62",
									 x"0AB42",x"0A342",x"10000",x"0A322",x"09B22",x"09B02",x"09AE2",x"08AC1",x"082A1",x"07A40",
									 x"08281",x"09BA4",x"0DDC7",x"0F6C7",x"0FEE7",x"0FE87",x"0FE47",x"0FE67",x"0FE47",x"1001B",
									 x"0FE67",x"0FEC8",x"10000",x"0E5E7",x"0ABE4",x"07A82",x"07A41",x"08281",x"092C1",x"092C2",
									 x"09B02",x"0A322",x"10000",x"0A342",x"0AB42",x"10000",x"0AB62",x"10000",x"0A342",x"10001",
									 x"0A322",x"09B02",x"10000",x"092E2",x"08AC1",x"08281",x"07A41",x"082C2",x"0B465",x"0EE28",
									 x"0FEA8",x"0FE67",x"0FE47",x"10000",x"0FE67",x"10001",x"0FE48",x"0FE68",x"10003",x"0FE69",
									 x"10004",x"0FE89",x"10001",x"0FE8A",x"10002",x"0FE89",x"10008",x"0FE8A",x"0FE6A",x"10000",
									 x"0FE69",x"0FE68",x"0FE67",x"10000",x"0FE47",x"10004",x"0FE27",x"10000",x"0FE06",x"10001",
									 x"0FDE6",x"10000",x"0FDC6",x"10000",x"0FDA5",x"0FD85",x"0FD65",x"0FD44",x"0FD24",x"0FCE3",
									 x"0F4A3",x"0F443",x"0EC24",x"0ECA9",x"0E56F",x"0EEB7",x"0F79C",x"0F7BE",x"0FFDF",x"0FFFF",
									 x"10006",x"0FFFF",x"10007",x"0F7DF",x"0F7BE",x"0F75C",x"0EE97",x"0ED6F",x"0ECA8",x"0EC44",
									 x"0F442",x"0FCA3",x"0FCE4",x"0FD24",x"0FD44",x"0FD65",x"0FD85",x"0FDA5",x"0FDC6",x"10000",
									 x"0FDE6",x"0FE06",x"10000",x"0FE26",x"0FE27",x"10001",x"0FE47",x"10006",x"0FE68",x"0FE69",
									 x"10001",x"0FE89",x"10005",x"0FE8A",x"10001",x"0FE89",x"10001",x"0FE6A",x"10000",x"0FE89",
									 x"10002",x"0FE69",x"10000",x"0FE68",x"10005",x"0FE67",x"10000",x"0FE47",x"10003",x"0FE67",
									 x"0FEA8",x"0F688",x"0C526",x"09BA4",x"07A81",x"08281",x"08AA1",x"092C2",x"09AE2",x"09B02",
									 x"0A322",x"10000",x"0A342",x"0AB42",x"10000",x"0AB62",x"0AB42",x"0A342",x"10000",x"0A322",
									 x"09B22",x"09B02",x"092E1",x"08AC1",x"08281",x"07A60",x"08AE2",x"0AC24",x"0E608",x"0FEC8",
									 x"10000",x"0FE67",x"0FE47",x"1001D",x"0FE67",x"0FEA8",x"0FEC8",x"0EE28",x"0B465",x"082E2",
									 x"07A61",x"08281",x"092C1",x"092E1",x"09B02",x"09B22",x"0A322",x"0A342",x"10000",x"0AB42",
									 x"0AB62",x"10000",x"0A342",x"10001",x"0A322",x"09B02",x"10000",x"092E2",x"08AC1",x"08261",
									 x"07A61",x"09343",x"0C4E6",x"0F648",x"0FEA7",x"0FE46",x"0FE47",x"10000",x"0FE66",x"0FE67",
									 x"0FE47",x"10001",x"0FE68",x"10008",x"0FE89",x"10001",x"0FE8A",x"10003",x"0FE89",x"10008",
									 x"0FE6A",x"0FE69",x"0FE68",x"10000",x"0FE67",x"0FE47",x"10005",x"0FE27",x"10000",x"0FE26",
									 x"0FE06",x"10001",x"0FDE6",x"0FDC6",x"10000",x"0FDA5",x"0FD85",x"0FD65",x"0FD44",x"0FD24",
									 x"0FCE3",x"0F4A3",x"0F463",x"0F424",x"0ECA8",x"0E52D",x"0EE76",x"0F77C",x"0F7BE",x"0FFDF",
									 x"0FFFF",x"10006",x"0FFFF",x"10007",x"0F7DF",x"0F79E",x"0F73B",x"0EE55",x"0E50D",x"0EC87",
									 x"0EC44",x"0F462",x"0F4A3",x"0F4E3",x"0F524",x"0FD44",x"0FD64",x"0FD85",x"0FDA5",x"0FDC6",
									 x"10000",x"0FDE6",x"0FE06",x"10000",x"0FE26",x"0FE27",x"10001",x"0FE47",x"10005",x"0FE67",
									 x"0FE68",x"10002",x"0FE69",x"10003",x"0FE89",x"10004",x"0FE69",x"10003",x"0FE68",x"10004",
									 x"0FE67",x"10009",x"0FE47",x"0FE48",x"0FE67",x"0FEA8",x"0F6A8",x"0D586",x"0AC45",x"07A81",
									 x"07A41",x"08A82",x"092C2",x"092E2",x"09B22",x"0A322",x"10000",x"0A342",x"0AB42",x"10002",
									 x"0A342",x"10001",x"09B21",x"09B01",x"092E1",x"10000",x"07A60",x"07A80",x"09363",x"0B4A5",
									 x"0EE89",x"0FEA8",x"0FE87",x"0FE67",x"0FE47",x"1001C",x"0FE67",x"10000",x"0FEA8",x"0FEC8",
									 x"0F668",x"0BCE5",x"09363",x"07A81",x"07A41",x"08AC1",x"092E1",x"09B02",x"09B22",x"0A322",
									 x"0A342",x"0AB62",x"10001",x"0AB42",x"0AB62",x"10000",x"0A342",x"0A322",x"09B22",x"09B02",
									 x"092C1",x"08AA1",x"07A61",x"10000",x"0AC05",x"0D567",x"0F668",x"0FEA7",x"0FE46",x"0FE67",
									 x"10000",x"0FE66",x"0FE67",x"10001",x"0FE47",x"10000",x"0FE67",x"10003",x"0FE68",x"10000",
									 x"0FE67",x"0FE68",x"10000",x"0FE69",x"10007",x"0FE89",x"10002",x"0FE69",x"0FE89",x"10000",
									 x"0FE69",x"10000",x"0FE68",x"10000",x"0FE67",x"10000",x"0FE47",x"10006",x"0FE27",x"10000",
									 x"0FE26",x"0FE06",x"10000",x"0FDE6",x"0FDC6",x"0FDA5",x"10000",x"0FD85",x"0FD65",x"0FD44",
									 x"0FD24",x"0FCE4",x"0F4C3",x"0F483",x"0F444",x"0EC87",x"0ECEC",x"0EE14",x"0F73B",x"0F79D",
									 x"0F7BE",x"0FFFF",x"10006",x"0FFFF",x"10006",x"0FFDF",x"0F7DF",x"0F79E",x"0F71A",x"0EDF3",
									 x"0E4EB",x"0EC66",x"0F464",x"0F462",x"0F4A3",x"0F4E3",x"0F524",x"0FD64",x"0FD84",x"0FD85",
									 x"0FDA5",x"0FDC6",x"10000",x"0FDE6",x"0FE06",x"10000",x"0FE26",x"0FE27",x"10000",x"0FE47",
									 x"10007",x"0FE67",x"10001",x"0FE68",x"10000",x"0FE69",x"10003",x"0FE89",x"0FE69",x"10004",
									 x"0FE48",x"10000",x"0FE68",x"10000",x"0FE67",x"10003",x"0FE47",x"10007",x"0FE67",x"10000",
									 x"0FE47",x"0FE48",x"0FE67",x"0FE88",x"0FEA9",x"0E628",x"0CD27",x"082A1",x"07200",x"08261",
									 x"092E2",x"09B02",x"10001",x"0A342",x"0AB42",x"10000",x"0A342",x"0AB42",x"0AB62",x"0A362",
									 x"0A342",x"09B22",x"09B21",x"09B02",x"092E2",x"08AC2",x"07220",x"07A81",x"0A404",x"0CD45",
									 x"0FEC9",x"0FEA8",x"0FE67",x"0FE46",x"0FE47",x"1001C",x"0FE67",x"10000",x"0FE87",x"0FEA7",
									 x"0FEC9",x"0D5A7",x"0A404",x"07AA1",x"07221",x"08AA1",x"092E1",x"09B02",x"10000",x"09B22",
									 x"0A342",x"10000",x"0AB62",x"10000",x"0AB42",x"0A342",x"10001",x"09B22",x"09B01",x"09AE2",
									 x"092C2",x"08A81",x"07A21",x"07A81",x"0BCE6",x"0E628",x"0FEA8",x"10000",x"0FE67",x"0FE68",
									 x"0FE47",x"10006",x"0FE67",x"10000",x"0FE47",x"0FE67",x"10004",x"0FE68",x"10001",x"0FE69",
									 x"1000A",x"0FE68",x"10002",x"0FE67",x"10001",x"0FE47",x"10007",x"0FE27",x"10000",x"0FE06",
									 x"10000",x"0FDE6",x"0FDC6",x"0FDC5",x"0FDA5",x"0FD85",x"0FD65",x"0FD45",x"0FD44",x"0F504",
									 x"0F4C3",x"0F483",x"0F463",x"0F466",x"0ECCB",x"0EDD2",x"0F6FA",x"0F79D",x"0F7BE",x"0FFDF",
									 x"0FFFF",x"10005",x"0FFFF",x"10006",x"0FFDF",x"0F7BF",x"0F79E",x"0F6D9",x"0EDB1",x"0ECCA",
									 x"0EC66",x"0F464",x"0F483",x"0F4C3",x"0F504",x"0F524",x"0FD64",x"0FD84",x"0FD85",x"0FDA5",
									 x"0FDC6",x"10000",x"0FDE6",x"0FE06",x"10000",x"0FE26",x"0FE27",x"10001",x"0FE47",x"10006",
									 x"0FE67",x"10002",x"0FE68",x"1000F",x"0FE48",x"0FE47",x"1000E",x"0FE48",x"0FE47",x"0FE87",
									 x"0FEA8",x"0F6A9",x"0E5E9",x"08B01",x"07221",x"08261",x"08AC1",x"092E1",x"09B02",x"10000",
									 x"0A322",x"0A342",x"10002",x"0A362",x"0A342",x"09B22",x"10000",x"09B02",x"10000",x"092C2",
									 x"08AA2",x"07220",x"082E2",x"0B4C6",x"0DDE7",x"0FF09",x"0FEA8",x"0FE67",x"0FE46",x"0FE47",
									 x"1001C",x"0FE67",x"10001",x"0FE87",x"0FF0A",x"0DE28",x"0B4C5",x"08B03",x"071E1",x"08AA1",
									 x"092E0",x"09B22",x"09B02",x"09B22",x"0A342",x"10000",x"0A362",x"0A342",x"10002",x"0A322",
									 x"09B22",x"09B02",x"09AE2",x"092A2",x"08A62",x"07A41",x"082E2",x"0D5A8",x"0FECA",x"0FEA9",
									 x"0FE88",x"0FE68",x"0FE48",x"0FE47",x"10009",x"0FE67",x"10002",x"0FE47",x"0FE67",x"0FE47",
									 x"0FE67",x"10000",x"0FE68",x"1000C",x"0FE67",x"10003",x"0FE47",x"10008",x"0FE27",x"0FE26",
									 x"0FE06",x"10000",x"0FDE6",x"0FDC5",x"0FDA5",x"10000",x"0FD85",x"0FD65",x"0FD44",x"0F504",
									 x"0F4C3",x"0F4A3",x"0F463",x"0F445",x"0ECAA",x"0E571",x"0EED9",x"0F79D",x"0F7BE",x"0FFDF",
									 x"0FFFF",x"10005",x"0FFFF",x"10006",x"0FFDF",x"0F7BF",x"0EF9E",x"0EED9",x"0ED6F",x"0ECA9",
									 x"0EC45",x"0F463",x"0F483",x"0F4C3",x"0F504",x"0FD24",x"0FD64",x"0FD84",x"0FD85",x"0FDA5",
									 x"0FDC5",x"0FDC6",x"0FDE6",x"0FE06",x"10000",x"0FE26",x"0FE27",x"10000",x"0FE47",x"10008",
									 x"0FE67",x"10001",x"0FE47",x"0FE48",x"10001",x"0FE68",x"10004",x"0FE67",x"0FE47",x"10015",
									 x"0FE67",x"10000",x"0FE87",x"0FEA8",x"0FEEA",x"0EE4A",x"09BA3",x"07A81",x"07A61",x"08AA1",
									 x"092E1",x"09B01",x"10000",x"0A321",x"0A322",x"10001",x"0A342",x"10001",x"09B22",x"10001",
									 x"09B02",x"092C2",x"08281",x"07A41",x"09363",x"0C567",x"0E648",x"0FF09",x"0FEA8",x"0FE67",
									 x"0FE47",x"1001E",x"0FE48",x"0FE67",x"0FEA8",x"0FF0A",x"0E688",x"0CD66",x"09BA4",x"07A21",
									 x"08262",x"08AA0",x"09301",x"09B22",x"10001",x"0A342",x"10004",x"0A322",x"09B22",x"09302",
									 x"092E2",x"08AA1",x"08262",x"07A82",x"09362",x"0E628",x"0FEE9",x"0FEA9",x"0FE88",x"0FE48",
									 x"10001",x"0FE47",x"10010",x"0FE67",x"10002",x"0FE68",x"10005",x"0FE48",x"10000",x"0FE67",
									 x"0FE47",x"1000D",x"0FE27",x"10000",x"0FE06",x"10001",x"0FDE6",x"0FDC6",x"0FDA5",x"10000",
									 x"0FD85",x"0FD65",x"0FD45",x"0FD04",x"0FCE4",x"0F4A3",x"0F463",x"0EC64",x"0ECA9",x"0ED4F",
									 x"0EED8",x"0F79D",x"0F7BE",x"0FFDF",x"0FFFF",x"10005",x"0FFFF",x"10006",x"0FFDF",x"0F7BE",
									 x"0EF7E",x"0EEB8",x"0F52D",x"0ECA8",x"0EC45",x"0F463",x"0F4A3",x"0F4E4",x"0F504",x"0FD24",
									 x"0FD65",x"0FD85",x"0FDA5",x"10000",x"0FDC5",x"0FDC6",x"0FDE6",x"0FE06",x"10000",x"0FE26",
									 x"0FE27",x"10000",x"0FE47",x"1000F",x"0FE67",x"0FE47",x"1001B",x"0FE67",x"10001",x"0FEA8",
									 x"0FF09",x"0F6CA",x"0C526",x"09383",x"07240",x"07A40",x"092C2",x"09AE2",x"09AE1",x"09B01",
									 x"09B22",x"0A322",x"10002",x"09B22",x"10001",x"09B01",x"092E2",x"08260",x"07A60",x"082E1",
									 x"0AC65",x"0E669",x"0F6EA",x"0FF09",x"0FE87",x"0FE67",x"0FE47",x"10020",x"0FE88",x"0FEE9",
									 x"0FF09",x"0E689",x"0BCE6",x"082C2",x"07A40",x"08260",x"09301",x"10000",x"09B22",x"10001",
									 x"0A322",x"0A342",x"0A322",x"10001",x"09B21",x"09B01",x"092E1",x"092A1",x"08261",x"07240",
									 x"08B63",x"0BD06",x"0F6C9",x"0FF09",x"0FEC8",x"0FE88",x"0FE47",x"1001D",x"0FE67",x"0FE47",
									 x"10010",x"0FE27",x"10000",x"0FE06",x"10001",x"0FDE6",x"0FDC6",x"0FDA5",x"10000",x"0FD85",
									 x"0FD65",x"0FD45",x"0FD04",x"0FCE4",x"0F4A3",x"0F483",x"0EC64",x"0EC88",x"0E52E",x"0EEB7",
									 x"0F79D",x"0F79E",x"0FFDF",x"0FFFF",x"10005",x"0FFFF",x"10006",x"0FFDF",x"0F7BE",x"0EF7E",
									 x"0EE97",x"0ECEC",x"0EC67",x"0EC45",x"0F463",x"0F4C3",x"0F4E4",x"0FD24",x"0FD44",x"0FD65",
									 x"0FD85",x"0FDA5",x"10000",x"0FDC5",x"0FDC6",x"0FDE6",x"0FE06",x"10000",x"0FE26",x"0FE27",
									 x"10000",x"0FE47",x"1000F",x"0FE67",x"0FE47",x"1001C",x"0FE67",x"10000",x"0FE87",x"0FEC8",
									 x"0FF09",x"0EE89",x"0C507",x"09343",x"07A41",x"08241",x"09282",x"09AC2",x"09AE2",x"09B02",
									 x"09B01",x"09B02",x"09B22",x"10001",x"09B02",x"092E1",x"10000",x"08A81",x"08240",x"082C0",
									 x"0AC24",x"0DE08",x"0FF0A",x"0FF09",x"0FEA8",x"0FE67",x"0FE47",x"0FE67",x"0FE47",x"1001F",
									 x"0FE67",x"0FEA8",x"0FF09",x"0F72A",x"0DE28",x"0AC65",x"082C1",x"08260",x"08AA1",x"092C1",
									 x"092E1",x"09301",x"09B01",x"09B22",x"0A321",x"09B22",x"0A302",x"09B02",x"10000",x"09AE1",
									 x"092C1",x"08A61",x"08242",x"08B02",x"0BD06",x"0E669",x"0FF29",x"0FF08",x"0FE88",x"0FE67",
									 x"0FE47",x"1001D",x"0FE67",x"0FE47",x"10010",x"0FE27",x"10000",x"0FE06",x"10001",x"0FDE6",
									 x"0FDC6",x"0FDA5",x"10000",x"0FD85",x"10000",x"0FD65",x"0FD04",x"0FCE4",x"0F4C3",x"0F483",
									 x"0EC44",x"0EC66",x"0E4EC",x"0EE96",x"0F79D",x"0F79E",x"0FFDF",x"0FFFF",x"10005",x"0FFFF",
									 x"10006",x"0FFDF",x"0F7BE",x"0EF7D",x"0EE97",x"0E4CA",x"0EC46",x"0EC44",x"0F463",x"0F4C3",
									 x"0FCE4",x"0FD24",x"0FD44",x"0FD65",x"0FD85",x"0FDA5",x"0FDC5",x"10000",x"0FDE6",x"0FE06",
									 x"10001",x"0FE26",x"0FE27",x"10000",x"0FE47",x"10027",x"0FE67",x"10004",x"0FE47",x"10000",
									 x"0FE67",x"10000",x"0FEA8",x"0FF08",x"0FF2A",x"0E649",x"0BCC6",x"08AE2",x"079E0",x"08A41",
									 x"092A2",x"09AE2",x"09B02",x"09B01",x"09B02",x"09B22",x"09B02",x"10000",x"09302",x"092C1",
									 x"092C2",x"07A20",x"082A2",x"09B83",x"0CD87",x"0F6EA",x"0FF2A",x"0FEE8",x"0FE87",x"0FE67",
									 x"0FE47",x"0FE68",x"10000",x"0FE47",x"1001E",x"0FE67",x"0FE88",x"0FEE9",x"0FF29",x"0F72B",
									 x"0D5C9",x"09BC3",x"08AC1",x"07A00",x"08A81",x"092C1",x"092E1",x"09301",x"09B21",x"10001",
									 x"09B01",x"10000",x"09AE2",x"092C2",x"08A61",x"07A00",x"082A2",x"0B485",x"0DE28",x"0FF2A",
									 x"0FF28",x"0FEC8",x"0FE87",x"0FE47",x"10031",x"0FE27",x"10000",x"0FE06",x"10001",x"0FDE6",
									 x"0FDC6",x"0FDC5",x"0FDA5",x"0FD85",x"10000",x"0FD44",x"0FD24",x"0FCE4",x"0F4C3",x"0F483",
									 x"0EC44",x"0F445",x"0E4CA",x"0EE56",x"0F77D",x"0F79E",x"0FFDF",x"0FFFF",x"10005",x"0FFFF",
									 x"10006",x"0FFDF",x"0F7BE",x"0EF7D",x"0EE76",x"0ECA9",x"0EC45",x"0EC44",x"0F462",x"0F4C3",
									 x"0FCE4",x"0FD24",x"0FD44",x"0FD85",x"10000",x"0FDA5",x"0FDC5",x"10000",x"0FDE6",x"0FE06",
									 x"10001",x"0FE26",x"0FE27",x"10000",x"0FE47",x"10027",x"0FE67",x"10005",x"0FE47",x"10001",
									 x"0FE88",x"0FEE8",x"0FF49",x"0EEEA",x"0D5E8",x"0A403",x"07A80",x"08260",x"08241",x"08A81",
									 x"092C1",x"092E1",x"09B02",x"09B22",x"09302",x"092E2",x"08AA1",x"08260",x"08261",x"07A60",
									 x"09BA4",x"0BCE6",x"0E689",x"0FF2A",x"0FF09",x"0FEA8",x"0FE67",x"0FE47",x"10000",x"0FE48",
									 x"0FE47",x"10020",x"0FE87",x"0FEA8",x"0FF09",x"0FF4B",x"0E68A",x"0BD26",x"09BA3",x"07A40",
									 x"10000",x"08260",x"08AA1",x"092C1",x"09B02",x"10000",x"09B01",x"09B00",x"092C1",x"08AA1",
									 x"08261",x"07A40",x"082A1",x"09BC3",x"0CD87",x"0EEC9",x"0FF4A",x"0FEE8",x"0FEA8",x"0FE67",
									 x"0FE47",x"10001",x"0FE67",x"10000",x"0FE47",x"1002C",x"0FE27",x"10000",x"0FE26",x"0FE06",
									 x"10000",x"0FDE6",x"10000",x"0FDC6",x"0FDA5",x"0FD85",x"0FD84",x"0FD44",x"0FD24",x"0F504",
									 x"0F4C3",x"0F483",x"0F424",x"0F444",x"0E4C8",x"0EE35",x"0F77D",x"0F79E",x"0FFDF",x"0FFFF",
									 x"10005",x"0FFFF",x"10005",x"0FFDF",x"0F7BE",x"0F79E",x"0EF5D",x"0EE56",x"0EC88",x"0EC45",
									 x"0EC44",x"0F462",x"0F4C3",x"0FCE3",x"0FD24",x"0FD44",x"0FD84",x"0FD85",x"0FDA5",x"0FDC5",
									 x"10000",x"0FDE6",x"0FE06",x"10001",x"0FE26",x"0FE27",x"10000",x"0FE47",x"10027",x"0FE67",
									 x"10005",x"0FE47",x"10001",x"0FE68",x"0FEA8",x"0FF29",x"0FF4B",x"0FF2B",x"0DE29",x"0AC84",
									 x"09342",x"08261",x"10000",x"08A80",x"08AA1",x"08AC1",x"10001",x"08AA1",x"08281",x"07A81",
									 x"082C1",x"09BC3",x"0CDA8",x"0E6A9",x"0FF4A",x"10000",x"0FEC8",x"0FE88",x"0FE47",x"10001",
									 x"0FE68",x"0FE47",x"10020",x"0FE67",x"0FE87",x"0FEC7",x"0FF2A",x"0FF4B",x"0EEEA",x"0CDE8",
									 x"0A404",x"082A1",x"08260",x"08281",x"08A81",x"08AA1",x"092C2",x"092A1",x"10000",x"08AA1",
									 x"08260",x"07A80",x"08B21",x"0AC64",x"0D608",x"0F70B",x"0FF2A",x"0FF09",x"0FEA8",x"0FE67",
									 x"10000",x"0FE47",x"10002",x"0FE67",x"0FE47",x"1002C",x"0FE27",x"10000",x"0FE26",x"0FE06",
									 x"10000",x"0FDE6",x"10000",x"0FDC6",x"0FDC5",x"0FDA5",x"0FD85",x"0FD64",x"0FD24",x"0FD03",
									 x"0F4C3",x"0F483",x"0F424",x"0F423",x"0E4A7",x"0EE14",x"0F75D",x"0F79E",x"0FFDF",x"0FFFF",
									 x"10005",x"0FFFF",x"10006",x"0F7BE",x"0F79E",x"0EF5D",x"0EE35",x"0EC68",x"0EC24",x"0F444",
									 x"0F463",x"0F4C3",x"0FCE4",x"0FD24",x"0FD44",x"0FD84",x"0FD85",x"0FDA5",x"0FDC5",x"0FDC6",
									 x"0FDE6",x"0FE06",x"10001",x"0FE26",x"0FE27",x"10000",x"0FE47",x"10000",x"0FE48",x"10001",
									 x"0FE47",x"0FE48",x"0FE47",x"10023",x"0FE67",x"10000",x"0FE47",x"10004",x"0FE88",x"0FEC9",
									 x"0FF09",x"0FF4A",x"0FF6B",x"0E6AA",x"0CDA9",x"0B486",x"09BA4",x"08AE2",x"082A1",x"07A40",
									 x"07200",x"07A40",x"08AC1",x"09B63",x"0AC45",x"0B506",x"0D629",x"0F72B",x"0FF6A",x"0FF49",
									 x"0FF09",x"0FEA8",x"0FE67",x"0FE47",x"10001",x"0FE67",x"0FE47",x"1001F",x"0FE67",x"0FE47",
									 x"0FE67",x"0FEA7",x"0FEE8",x"0FF29",x"0FF6B",x"0F74B",x"0DE6A",x"0BD27",x"0AC45",x"09BA3",
									 x"082A1",x"07A41",x"07A01",x"10000",x"08262",x"08AE2",x"09383",x"0B4A5",x"0CDA8",x"0DE89",
									 x"0F74B",x"0FF6B",x"0FF29",x"0FEA8",x"0FE68",x"0FE47",x"10032",x"0FE27",x"10000",x"0FE26",
									 x"10000",x"0FE06",x"10000",x"0FDE6",x"10000",x"0FDC6",x"0FDC5",x"0FDA5",x"0FD85",x"0FD64",
									 x"0FD24",x"0FD04",x"0F4C3",x"0F483",x"0F423",x"10000",x"0EC66",x"0EDF3",x"0EF5C",x"0EF9E",
									 x"0F7BE",x"0FFDF",x"0FFFF",x"10004",x"0FFFF",x"10006",x"0F7BE",x"0F79E",x"0E75C",x"0EE34",
									 x"0EC67",x"0F424",x"0F444",x"0F463",x"0F4C3",x"0FCE4",x"0FD24",x"0FD44",x"0FD84",x"0FD85",
									 x"0FDA5",x"0FDC6",x"10000",x"0FDE6",x"0FE06",x"10001",x"0FE26",x"0FE27",x"10000",x"0FE47",
									 x"10032",x"0FE67",x"0FE87",x"0FEC8",x"0FF29",x"0FF8B",x"0FF8C",x"0EF2B",x"0D649",x"0B506",
									 x"09BC3",x"08B21",x"07AC0",x"07A80",x"082E1",x"09382",x"0AC84",x"0CDC7",x"0DE89",x"0F76C",
									 x"0FFAB",x"0FF6A",x"0FF09",x"0FEA8",x"0FE87",x"0FE67",x"0FE47",x"10026",x"0FE67",x"0FE87",
									 x"0FF09",x"0FF4A",x"0FF8C",x"10000",x"0DEA9",x"0CDE7",x"0B4E5",x"09382",x"082E1",x"07A60",
									 x"07AA1",x"08322",x"093C3",x"0ACA5",x"0D608",x"0EF0A",x"0FF8B",x"0FF8A",x"0FF49",x"0FEC8",
									 x"0FE67",x"0FE47",x"10033",x"0FE27",x"10000",x"0FE26",x"10000",x"0FE06",x"10000",x"0FDE6",
									 x"10000",x"0FDC6",x"0FDC5",x"0FDA5",x"0FD85",x"0FD44",x"0FD24",x"0FD04",x"0F4C3",x"0FC83",
									 x"0F443",x"0F442",x"0F446",x"0EDF3",x"0EF5C",x"0EF7D",x"0F7BE",x"0FFDF",x"0FFFF",x"10004",
									 x"0FFFF",x"10005",x"0FFDF",x"0F7BE",x"0F79E",x"0E75C",x"0EE34",x"0EC67",x"0F423",x"0F444",
									 x"0F483",x"0F4C3",x"0FCE4",x"0FD24",x"0FD44",x"0FD84",x"0FD85",x"0FDA5",x"0FDC6",x"10000",
									 x"0FDE6",x"0FE06",x"10001",x"0FE26",x"0FE27",x"10000",x"0FE47",x"10033",x"0FE67",x"0FEA8",
									 x"0FEE8",x"0FF29",x"0FF8A",x"0FF8B",x"0F76B",x"0E6EA",x"0DEAA",x"0DE69",x"0D629",x"10001",
									 x"0DE69",x"0EF0A",x"0F76B",x"10000",x"0FF8B",x"0FF6A",x"0FF09",x"0FEC8",x"0FE68",x"0FE67",
									 x"0FE47",x"10028",x"0FE68",x"0FEC8",x"0FEE9",x"0FF4A",x"0FF8B",x"10000",x"0F74A",x"0EEEA",
									 x"0DE89",x"0DE49",x"0D629",x"10000",x"0DE6A",x"0DE8A",x"0E6CA",x"0F74A",x"0FF8A",x"10000",
									 x"0FF49",x"0FEE9",x"0FE88",x"0FE47",x"10034",x"0FE27",x"10000",x"0FE26",x"10000",x"0FE06",
									 x"10000",x"0FDE6",x"10000",x"0FDC6",x"0FDC5",x"0FDA5",x"0FD85",x"0FD44",x"0FD24",x"0FD04",
									 x"0F4E3",x"0FC83",x"0F443",x"0F442",x"0F426",x"0EDD2",x"0EF5C",x"0EF7D",x"0F7BE",x"0FFDF",
									 x"0FFFF",x"10004",x"0FFFF",x"10005",x"0FFDF",x"0F7BE",x"0EF7D",x"0E75C",x"0EE34",x"0EC46",
									 x"0F423",x"0F443",x"0F483",x"0F4C3",x"0FD04",x"0FD24",x"0FD44",x"0FD84",x"0FD85",x"0FDA5",
									 x"0FDC6",x"10000",x"0FE06",x"10002",x"0FE26",x"0FE27",x"10000",x"0FE47",x"10003",x"0FE27",
									 x"0FE47",x"1002D",x"0FE67",x"0FE87",x"0FEA8",x"0FEC8",x"0FF09",x"0FF49",x"0FFAB",x"0FFCB",
									 x"0FFCC",x"10005",x"0FFAB",x"0FF8A",x"0FF29",x"0FEE8",x"0FEC8",x"0FE88",x"0FE47",x"10000",
									 x"0FE67",x"0FE47",x"10000",x"0FE67",x"10000",x"0FE47",x"10022",x"0FE48",x"10000",x"0FE88",
									 x"0FEA8",x"0FEC8",x"0FF09",x"0FF8A",x"0FF8B",x"0FFAB",x"0FFCC",x"10000",x"0FFCD",x"0FFCC",
									 x"0FFCD",x"0FFCC",x"0FFAC",x"0FF8B",x"0FF4A",x"0FF29",x"0FEC8",x"0FEA8",x"0FE67",x"0FE47",
									 x"10034",x"0FE27",x"10001",x"0FE26",x"0FE06",x"10000",x"0FDE6",x"0FDC6",x"10000",x"0FDA5",
									 x"0FD85",x"0FD84",x"0FD44",x"0FD24",x"0FD04",x"0F4E3",x"0FC83",x"0F443",x"0F422",x"0F425",
									 x"0EDD2",x"0EF5C",x"0EF7D",x"0F7BE",x"0FFDF",x"0FFFF",x"10004",x"0FFFF",x"10005",x"0FFDF",
									 x"0F7BE",x"0EF7D",x"0E75C",x"0EE33",x"0EC25",x"0F422",x"0F443",x"0F483",x"0F4C3",x"0FD04",
									 x"0FD24",x"0FD44",x"0FD84",x"0FD85",x"0FDA5",x"0FDC6",x"10000",x"0FDE6",x"0FE06",x"10001",
									 x"0FE26",x"0FE27",x"10001",x"0FE47",x"10034",x"0FE67",x"0FE88",x"0FEA9",x"0FEE9",x"0FF2A",
									 x"0FF4A",x"0FF8B",x"10000",x"0FFAB",x"10001",x"0FF8B",x"0FF6B",x"0FF4A",x"0FF09",x"0FEE8",
									 x"0FEA8",x"0FE87",x"0FE67",x"0FE47",x"10002",x"0FE67",x"10001",x"0FE47",x"10022",x"0FE48",
									 x"10000",x"0FE67",x"0FE87",x"0FEA8",x"0FEC8",x"0FF09",x"0FF2A",x"0FF6B",x"0FF8B",x"0FFAB",
									 x"0FFAC",x"0FFAB",x"10000",x"0FF8B",x"0FF6B",x"0FF2A",x"0FEE9",x"0FEC8",x"0FE88",x"0FE67",
									 x"10000",x"0FE47",x"10035",x"0FE27",x"10001",x"0FE06",x"10000",x"0FDE6",x"0FDC6",x"0FDC5",
									 x"0FDA5",x"10000",x"0FD64",x"0FD44",x"0FD24",x"0FD04",x"0F4E3",x"0F4A3",x"0F443",x"0F422",
									 x"0F425",x"0EDD2",x"0EF5C",x"0EF7D",x"0F7BE",x"0FFDF",x"0FFFF",x"10004",x"0FFFF",x"10005",
									 x"0FFDF",x"0F7BE",x"0EF7E",x"0E75C",x"0EE13",x"0EC24",x"0F422",x"0F463",x"0F483",x"0F4C3",
									 x"0FD04",x"0FD24",x"0FD44",x"0FD84",x"0FD85",x"0FDA5",x"0FDC6",x"10000",x"0FDE6",x"0FE06",
									 x"10001",x"0FE26",x"0FE27",x"10001",x"0FE47",x"10035",x"0FE67",x"0FE68",x"0FE88",x"0FEC8",
									 x"0FEE9",x"0FF09",x"10000",x"0FF2A",x"10000",x"0FF29",x"10000",x"0FEE9",x"0FEC9",x"0FEA9",
									 x"0FE88",x"0FE67",x"10001",x"0FE47",x"10001",x"0FE67",x"10002",x"0FE47",x"10024",x"0FE67",
									 x"10000",x"0FE87",x"0FE88",x"0FEA8",x"0FEC9",x"0FEE9",x"0FF0A",x"0FF2A",x"0FF4A",x"10000",
									 x"0FF2A",x"0FF09",x"0FEE9",x"0FEC8",x"0FEA8",x"0FE87",x"0FE47",x"10038",x"0FE27",x"10001",
									 x"0FE06",x"10000",x"0FDE6",x"0FDC6",x"0FDC5",x"0FDA5",x"10000",x"0FD64",x"10000",x"0FD24",
									 x"0FD04",x"0F4E3",x"0F4A3",x"0F463",x"0F422",x"0F425",x"0F5B2",x"0EF5C",x"0EF7D",x"0F7BE",
									 x"0FFDF",x"0FFFF",x"10004",x"0FFFF",x"10005",x"0FFDF",x"0F7BE",x"0EF7E",x"0EF5C",x"0EE13",
									 x"0EC24",x"0F402",x"0F443",x"0F483",x"0F4C3",x"0FD04",x"0FD24",x"0FD44",x"0FD84",x"0FD85",
									 x"0FDA5",x"0FDC6",x"10000",x"0FDE6",x"0FE06",x"10001",x"0FE26",x"0FE27",x"10001",x"0FE47",
									 x"10037",x"0FE67",x"10000",x"0FE87",x"10000",x"0FE88",x"0FEA8",x"10000",x"0FEA7",x"10000",
									 x"0FE87",x"0FE67",x"0FE48",x"0FE47",x"10006",x"0FE67",x"10001",x"0FE47",x"10024",x"0FE67",
									 x"10001",x"0FE47",x"0FE67",x"10000",x"0FE88",x"10001",x"0FEA8",x"10000",x"0FEA7",x"0FE87",
									 x"10000",x"0FE67",x"10000",x"0FE47",x"0FE27",x"0FE47",x"1001C",x"0FE27",x"0FE47",x"10014",
									 x"0FE27",x"10005",x"0FE06",x"10000",x"0FDE6",x"0FDC6",x"10000",x"0FDA5",x"10000",x"0FD65",
									 x"0FD64",x"0FD24",x"0FD04",x"0F4E3",x"0F4A3",x"0F463",x"0F422",x"0F424",x"0EDB1",x"0EF5C",
									 x"0EF7E",x"0F7BE",x"0FFDF",x"0FFFF",x"10004",x"0FFFF",x"10005",x"0FFDF",x"0F7BE",x"0EF7E",
									 x"0EF3C",x"0EE13",x"0EC24",x"0F402",x"0F443",x"0F483",x"0F4C3",x"0FD04",x"0FD24",x"0FD44",
									 x"0FD84",x"0FD85",x"0FDA5",x"0FDC5",x"0FDC6",x"0FDE6",x"0FE06",x"10001",x"0FE26",x"0FE27",
									 x"10001",x"0FE47",x"1003A",x"0FE67",x"10004",x"0FE47",x"1000C",x"0FE67",x"1001C",x"0FE47",
									 x"1000D",x"0FE67",x"10004",x"0FE47",x"1001D",x"0FE27",x"10004",x"0FE47",x"10012",x"0FE27",
									 x"10004",x"0FE06",x"0FE27",x"0FE07",x"0FE06",x"0FDE6",x"10000",x"0FDC6",x"0FDC5",x"0FDA5",
									 x"0FD85",x"0FD65",x"0FD24",x"0FD04",x"0F4E4",x"0FCA3",x"0F442",x"0EC22",x"0EC24",x"0EDD0",
									 x"0EF3C",x"0EF7E",x"0F7BE",x"0FFDF",x"0FFFF",x"10004",x"0FFFF",x"10005",x"0FFDF",x"0F7BE",
									 x"0EF7E",x"0E73C",x"0EE12",x"0EC04",x"0F402",x"0F443",x"0F483",x"0F4C3",x"0FD04",x"0FD24",
									 x"0FD44",x"0FD84",x"0FD85",x"0FDA5",x"0FDC5",x"0FDC6",x"0FDE6",x"0FE06",x"10001",x"0FE26",
									 x"0FE27",x"10001",x"0FE47",x"1003B",x"0FE67",x"10001",x"0FE47",x"1000D",x"0FE67",x"1001E",
									 x"0FE47",x"10009",x"0FE67",x"0FE47",x"10002",x"0FE67",x"10000",x"0FE47",x"1002B",x"0FE27",
									 x"10001",x"0FE47",x"10007",x"0FE27",x"10006",x"0FE06",x"0FE26",x"0FE06",x"10000",x"0FDE6",
									 x"10000",x"0FDC6",x"0FDC5",x"0FDA5",x"0FD85",x"0FD44",x"0FD24",x"0FD04",x"0F4E4",x"0FCA3",
									 x"0F462",x"0F422",x"0EC04",x"0EDD0",x"0EF3C",x"0EF7E",x"0F7BE",x"0FFDF",x"0FFFF",x"10004",
									 x"0FFFF",x"10005",x"0FFDF",x"0F7BE",x"0EF7E",x"0E73C",x"0EE12",x"0EC04",x"0F402",x"0F443",
									 x"0F483",x"0F4E3",x"0FD04",x"0FD24",x"0FD44",x"0FD84",x"0FD85",x"0FDA5",x"0FDC5",x"0FDC6",
									 x"0FDE6",x"0FE06",x"10001",x"0FE26",x"0FE27",x"10001",x"0FE47",x"0FE27",x"10004",x"0FE47",
									 x"10032",x"0FE67",x"10001",x"0FE47",x"10000",x"0FE67",x"0FE47",x"1000C",x"0FE67",x"1001E",
									 x"0FE47",x"1000B",x"0FE67",x"0FE47",x"10000",x"0FE67",x"0FE47",x"10002",x"0FE67",x"10002",
									 x"0FE47",x"1000A",x"0FE27",x"10000",x"0FE47",x"10016",x"0FE27",x"10012",x"0FE06",x"0FE26",
									 x"0FE06",x"10000",x"0FDE6",x"10000",x"0FDC6",x"0FDA5",x"10000",x"0FD85",x"0FD44",x"0FD24",
									 x"0F504",x"0F4C4",x"0F4A3",x"0F462",x"0F422",x"0EC24",x"0F5D0",x"0EF3C",x"0EF7E",x"0F7BE",
									 x"0FFDF",x"0FFFF",x"10004",x"0FFFF",x"10005",x"0FFDF",x"0F7BE",x"0EF7D",x"0E73C",x"0EE12",
									 x"0EC24",x"0F401",x"0F443",x"0F483",x"0FCE4",x"0FD04",x"0FD24",x"0FD44",x"0FD84",x"0FD85",
									 x"0FDA5",x"0FDC6",x"10000",x"0FDE6",x"0FE06",x"10001",x"0FE26",x"0FE27",x"10008",x"0FE47",
									 x"10033",x"0FE67",x"10000",x"0FE47",x"1000F",x"0FE67",x"10030",x"0FE47",x"1002B",x"0FE27",
									 x"10011",x"0FE06",x"10003",x"0FDE6",x"10001",x"0FDA5",x"10000",x"0FD65",x"0FD44",x"0FD24",
									 x"0FD04",x"0F4E4",x"0F4A3",x"0F462",x"0EC22",x"0EC04",x"0EDD0",x"0EF3C",x"0EF7E",x"0F7BE",
									 x"0FFDF",x"0FFFF",x"10004",x"0FFFF",x"10005",x"0FFDF",x"0F7BE",x"0EF7D",x"0E73C",x"0EE12",
									 x"0EC24",x"0F401",x"0F443",x"0F483",x"0F4C3",x"0FCE4",x"0FD24",x"0FD44",x"0FD64",x"0FD85",
									 x"0FDA5",x"10000",x"0FDC6",x"0FDE6",x"0FE06",x"10002",x"0FE26",x"0FE27",x"1000D",x"0FE47",
									 x"10004",x"0FE27",x"10001",x"0FE47",x"10008",x"0FE46",x"10001",x"0FE47",x"10017",x"0FE67",
									 x"10000",x"0FE47",x"1000F",x"0FE67",x"1002A",x"0FE47",x"10017",x"0FE46",x"10001",x"0FE47",
									 x"10004",x"0FE46",x"10009",x"0FE26",x"10001",x"0FE27",x"10014",x"0FE06",x"10003",x"0FDE6",
									 x"0FDE5",x"0FDC5",x"0FDA5",x"10000",x"0FD85",x"0FD44",x"0FD24",x"0FD04",x"0F4E4",x"0F4A3",
									 x"0F462",x"0F422",x"0EC04",x"0EDB0",x"0EF3C",x"0EF7E",x"0F7BE",x"0FFDF",x"0FFFF",x"10004",
									 x"0FFFF",x"10005",x"0FFDF",x"0F7BE",x"0EF7E",x"0E73C",x"0EE13",x"0EC24",x"0F402",x"0F463",
									 x"0F483",x"0F4C3",x"0F4E4",x"0FD24",x"0FD44",x"0FD64",x"0FD84",x"0FDA5",x"10000",x"0FDC5",
									 x"0FDE6",x"0FE06",x"10002",x"0FE26",x"10000",x"0FE27",x"1000C",x"0FE47",x"10003",x"0FE27",
									 x"10000",x"0FE26",x"10000",x"0FE27",x"0FE47",x"10006",x"0FE26",x"0FE46",x"10001",x"0FE47",
									 x"1001F",x"0FE46",x"10003",x"0FE47",x"10004",x"0FE67",x"1001E",x"0FE66",x"1000A",x"0FE46",
									 x"10003",x"0FE47",x"10005",x"0FE46",x"10003",x"0FE47",x"10006",x"0FE46",x"10001",x"0FE47",
									 x"10004",x"0FE46",x"10009",x"0FE26",x"10001",x"0FE27",x"10013",x"0FE26",x"0FE06",x"10003",
									 x"0FDE6",x"0FDC5",x"10000",x"0FDA5",x"0FD85",x"0FD65",x"0FD44",x"0FD24",x"0FD04",x"0F4E3",
									 x"0F4A3",x"0F442",x"0F422",x"0EC24",x"0EDD0",x"0EF3C",x"0EF5E",x"0F79E",x"0FFDF",x"0FFFF",
									 x"10004",x"0FFFF",x"10005",x"0FFDF",x"0F7BE",x"0EF7E",x"0E73C",x"0EE13",x"0EC45",x"0F422",
									 x"0F463",x"0F4A3",x"0F4C4",x"0F4E4",x"0FD24",x"0FD44",x"0FD84",x"0FD85",x"0FDA5",x"10000",
									 x"0FDC5",x"0FDE5",x"0FDE6",x"0FE06",x"10001",x"0FE26",x"10008",x"0FE27",x"1000A",x"0FE26",
									 x"10003",x"0FE46",x"0FE47",x"10002",x"0FE26",x"10003",x"0FE46",x"0FE47",x"10012",x"0FE46",
									 x"10001",x"0FE47",x"10007",x"0FE67",x"10036",x"0FE46",x"10003",x"0FE47",x"10011",x"0FE46",
									 x"0FE26",x"0FE46",x"0FE47",x"10004",x"0FE46",x"10004",x"0FE47",x"10004",x"0FE26",x"10007",
									 x"0FE27",x"10004",x"0FE26",x"10008",x"0FE06",x"10003",x"0FDE6",x"0FDC5",x"10000",x"0FDA5",
									 x"0FD84",x"0FD64",x"0FD44",x"0FD04",x"10000",x"0F4E3",x"0F483",x"0F443",x"0F441",x"0EC45",
									 x"0EDD1",x"0EF3B",x"0EF5D",x"0F79E",x"0FFDF",x"0FFFF",x"10004",x"0FFFF",x"10005",x"0FFDF",
									 x"0F7BE",x"0EF7D",x"0E73C",x"0EE13",x"0EC66",x"0F423",x"0F463",x"0F483",x"0F4C3",x"0FCE4",
									 x"0FD24",x"0FD44",x"0FD84",x"0FD85",x"0FDA5",x"10000",x"0FDC5",x"0FDE5",x"0FDE6",x"0FE06",
									 x"10001",x"0FE26",x"10019",x"0FE46",x"10003",x"0FE26",x"0FE46",x"10003",x"0FE47",x"10012",
									 x"0FE46",x"0FE66",x"0FE46",x"0FE47",x"10058",x"0FE46",x"10000",x"0FE47",x"10003",x"0FE46",
									 x"1000B",x"0FE26",x"10017",x"0FE06",x"10002",x"0FDE6",x"0FDE5",x"0FDC5",x"10000",x"0FDA5",
									 x"0FD84",x"0FD64",x"0FD44",x"0FD04",x"10000",x"0F4E3",x"0F483",x"0F443",x"0EC42",x"0EC45",
									 x"0EDD2",x"0EF3B",x"0EF5D",x"0F7BE",x"0FFDF",x"0FFFF",x"10004",x"0FFFF",x"10005",x"0FFDF",
									 x"0F7BE",x"0EF7D",x"0E73C",x"0E614",x"0EC67",x"0EC23",x"0F463",x"0F483",x"0F4C3",x"0FCE3",
									 x"0FD24",x"0FD44",x"0FD84",x"10000",x"0FDA5",x"10000",x"0FDC5",x"0FDE5",x"0FDE6",x"0FE06",
									 x"10001",x"0FE26",x"10019",x"0FE46",x"0FE26",x"10003",x"0FE46",x"10023",x"0FE47",x"1003C",
									 x"0FE46",x"10022",x"0FE26",x"1001B",x"0FE06",x"10001",x"0FDE6",x"0FDE5",x"0FDC5",x"10000",
									 x"0FDA5",x"0FD84",x"0FD64",x"0FD44",x"0FD24",x"0FD04",x"0F4E3",x"0F483",x"0F443",x"0EC42",
									 x"0EC66",x"0EDD2",x"0EF3B",x"0EF5D",x"0F7BE",x"0FFFF",x"10005",x"0FFFF",x"10006",x"0F7BE",
									 x"0EF7D",x"0E73C",x"0E614",x"0EC68",x"0EC24",x"0F464",x"0F482",x"0F4C3",x"0F4E3",x"0FD23",
									 x"0FD44",x"0FD84",x"10000",x"0FDA5",x"10000",x"0FDC5",x"10000",x"0FDE6",x"0FE06",x"10001",
									 x"0FE26",x"1001A",x"0FE46",x"1001F",x"0FE66",x"0FE46",x"10003",x"0FE66",x"10038",x"0FE46",
									 x"0FE47",x"10003",x"0FE66",x"10002",x"0FE46",x"10000",x"0FE66",x"10003",x"0FE46",x"10018",
									 x"0FE26",x"1001B",x"0FE06",x"10001",x"0FDE6",x"0FDC5",x"10000",x"0FDA5",x"10000",x"0FD84",
									 x"0FD64",x"0FD44",x"0FD24",x"0FD04",x"0F4E3",x"0FC84",x"0F443",x"0EC43",x"0EC66",x"0EDD3",
									 x"0EF3C",x"0EF7D",x"0F7BE",x"0FFFF",x"10005",x"0FFFF",x"10006",x"0F7BE",x"0EF7D",x"0E71B",
									 x"0E615",x"0EC88",x"0EC45",x"0F464",x"0F482",x"0F4C3",x"0F4E3",x"0FD23",x"0FD43",x"0FD64",
									 x"0FD84",x"0FD85",x"0FDA5",x"0FDC5",x"10000",x"0FDE6",x"0FE06",x"10002",x"0FE26",x"10019",
									 x"0FE46",x"10019",x"0FE66",x"10002",x"0FE46",x"0FE66",x"10049",x"0FE46",x"0FE66",x"10004",
									 x"0FE46",x"10018",x"0FE26",x"1001A",x"0FE06",x"10002",x"0FDE6",x"0FDC5",x"0FDA5",x"10001",
									 x"0FD84",x"0FD64",x"0FD44",x"0FD24",x"0FD04",x"0F4C3",x"0F464",x"0F444",x"0EC63",x"0EC67",
									 x"0EDD3",x"0EF3C",x"0EF7D",x"0F7BE",x"0FFFF",x"10005",x"0FFFF",x"10006",x"0F7BE",x"0EF7D",
									 x"0E71B",x"0E635",x"0E489",x"0EC45",x"0F464",x"0F483",x"0F4C3",x"0F4E3",x"0FD23",x"0FD44",
									 x"0FD64",x"0FD84",x"0FD85",x"0FDA5",x"10000",x"0FDC5",x"0FDE6",x"10000",x"0FE06",x"10001",
									 x"0FE26",x"10007",x"0FE46",x"10009",x"0FE26",x"10001",x"0FE46",x"1001D",x"0FE66",x"10002",
									 x"0FE46",x"0FE66",x"1000D",x"0FE65",x"0FE66",x"10039",x"0FE46",x"0FE66",x"10005",x"0FE46",
									 x"1001A",x"0FE26",x"0FE46",x"0FE26",x"10015",x"0FE06",x"10001",x"0FDE6",x"10000",x"0FDC5",
									 x"0FDA5",x"10001",x"0FD84",x"0FD64",x"0FD44",x"0FD24",x"0FD04",x"0F4C3",x"0F484",x"0F444",
									 x"0EC64",x"0E488",x"0EDD4",x"0EF3C",x"0EF7D",x"0F7BE",x"0FFFF",x"10005",x"0FFFF",x"10005",
									 x"0FFDF",x"0F7BE",x"0EF7D",x"0EF1B",x"0E635",x"0DCAA",x"0EC45",x"0F443",x"0F483",x"0F4C3",
									 x"0FCE3",x"0FD23",x"0FD44",x"0FD64",x"0FD84",x"0FD85",x"0FDA5",x"0FDC5",x"10000",x"0FDE5",
									 x"0FE05",x"10002",x"0FE26",x"10004",x"0FE46",x"1000B",x"0FE26",x"0FE47",x"10001",x"0FE46",
									 x"10004",x"0FE26",x"10000",x"0FE46",x"0FE45",x"0FE46",x"1000A",x"0FE66",x"0FE46",x"10008",
									 x"0FE66",x"1000F",x"0FE65",x"10001",x"0FE66",x"10034",x"0FE65",x"10001",x"0FE66",x"10008",
									 x"0FE46",x"10006",x"0FE66",x"10001",x"0FE46",x"10009",x"0FE45",x"0FE46",x"10002",x"0FE45",
									 x"0FE46",x"10000",x"0FE26",x"0FE46",x"0FE26",x"10012",x"0FE06",x"10002",x"0FDE5",x"0FDC5",
									 x"10000",x"0FDA5",x"0FD85",x"0FD84",x"0FD64",x"0FD44",x"0FD23",x"0FCE3",x"0FCC3",x"0F483",
									 x"0F443",x"0EC45",x"0DCA9",x"0E614",x"0EF3B",x"0EF5D",x"0F7BE",x"0FFFF",x"10005",x"0FFFF",
									 x"10006",x"0F7BE",x"0EF7D",x"0E71B",x"0E655",x"0E4EB",x"0EC66",x"0EC44",x"0F483",x"0F4A3",
									 x"0FCE3",x"0FD03",x"0FD43",x"0FD64",x"0FD84",x"0FD85",x"0FDA5",x"10000",x"0FDC5",x"0FDE5",
									 x"10000",x"0FE05",x"10000",x"0FE25",x"10000",x"0FE26",x"10002",x"0FE46",x"10002",x"0FE26",
									 x"10007",x"0FE46",x"10002",x"0FE47",x"10000",x"0FE46",x"10006",x"0FE26",x"0FE25",x"0FE46",
									 x"1000D",x"0FE66",x"10004",x"0FE46",x"0FE66",x"10008",x"0FE86",x"0FE66",x"10004",x"0FE86",
									 x"0FE85",x"10000",x"0FE86",x"10000",x"0FE65",x"1001B",x"0FE85",x"1000A",x"0FE65",x"10003",
									 x"0FE66",x"10002",x"0FE86",x"0FE66",x"0FE65",x"10002",x"0FE66",x"10012",x"0FE46",x"10000",
									 x"0FE45",x"10000",x"0FE46",x"0FE45",x"0FE26",x"10000",x"0FE46",x"10001",x"0FE45",x"10000",
									 x"0FE46",x"10002",x"0FE26",x"0FE46",x"0FE45",x"0FE46",x"0FE26",x"10012",x"0FE06",x"10001",
									 x"0FDE6",x"0FDE5",x"0FDC5",x"10000",x"0FDA5",x"0FD85",x"0FD64",x"10000",x"0FD43",x"0FD03",
									 x"0FCE3",x"0F4C3",x"0F483",x"0F443",x"0EC45",x"0E4CA",x"0E634",x"0E73B",x"0EF5D",x"0F7BE",
									 x"0FFFF",x"10005",x"0FFFF",x"10006",x"0FFDF",x"0EF7D",x"0E73B",x"0E656",x"0E50D",x"0EC87",
									 x"0EC44",x"0F483",x"0FCA3",x"0FCE3",x"0FD03",x"0FD23",x"0FD64",x"10000",x"0FD84",x"0FDA5",
									 x"10000",x"0FDC5",x"0FDE5",x"10000",x"0FE05",x"10000",x"0FE25",x"10001",x"0FE26",x"10001",
									 x"0FE46",x"10002",x"0FE26",x"10006",x"0FE25",x"0FE45",x"0FE25",x"0FE24",x"10000",x"0FE45",
									 x"0FE46",x"10000",x"0FE66",x"0FE65",x"0FE45",x"10001",x"0FE46",x"0FE45",x"10000",x"0FE25",
									 x"0FE45",x"0FE46",x"0FE45",x"10001",x"0FE46",x"10008",x"0FE66",x"10004",x"0FE46",x"0FE66",
									 x"10008",x"0FE86",x"0FE66",x"10003",x"0FE86",x"0FE85",x"10003",x"0FE86",x"0FE65",x"10019",
									 x"0FE85",x"1000B",x"0FE65",x"10003",x"0FE66",x"10002",x"0FE86",x"0FE66",x"0FE65",x"10003",
									 x"0FE66",x"10012",x"0FE65",x"10000",x"0FE45",x"10002",x"0FE25",x"0FE45",x"0FE65",x"10004",
									 x"0FE66",x"0FE45",x"10003",x"0FE25",x"0FE45",x"0FE46",x"0FE26",x"1000C",x"0FE25",x"0FE26",
									 x"10000",x"0FE05",x"10001",x"0FDE5",x"0FDC5",x"10001",x"0FDA5",x"0FD85",x"0FD64",x"10000",
									 x"0FD43",x"0FD03",x"0FCE3",x"0F4A3",x"0F483",x"0EC44",x"0EC66",x"0E4EB",x"0E634",x"0E73B",
									 x"0EF7D",x"0F7BE",x"0FFFF",x"10005",x"0FFFF",x"10006",x"0FFDF",x"0EF9D",x"0E73C",x"0E677",
									 x"0E52E",x"0EC88",x"0EC45",x"0F483",x"0FCA3",x"0FCC3",x"0FD03",x"0FD24",x"0FD64",x"0FD84",
									 x"10000",x"0FDA5",x"10000",x"0FDC4",x"0FDE5",x"10000",x"0FE05",x"10000",x"0FE25",x"0FE26",
									 x"0FE05",x"0FE26",x"0FE46",x"10001",x"0FE26",x"10000",x"0FE46",x"0FE26",x"10005",x"0FE25",
									 x"0FE45",x"10002",x"0FE65",x"0FE44",x"0FE25",x"0FE26",x"0FE46",x"0FE45",x"0FE66",x"10000",
									 x"0FE86",x"0FE85",x"10000",x"0FE65",x"10002",x"0FE45",x"10001",x"0FE65",x"10002",x"0FE45",
									 x"10000",x"0FE65",x"10020",x"0FE85",x"10026",x"0FE65",x"1001E",x"0FE66",x"0FE65",x"0FE45",
									 x"10001",x"0FE65",x"10004",x"0FE85",x"10001",x"0FE86",x"0FE66",x"0FE65",x"0F645",x"0F646",
									 x"0FE46",x"0FE65",x"10000",x"0FE45",x"10001",x"0FE25",x"10004",x"0FE26",x"10003",x"0FE25",
									 x"10005",x"0FE05",x"10001",x"0FDE5",x"10001",x"0FDC5",x"10000",x"0FDA5",x"0FD84",x"0FD64",
									 x"10000",x"0FD43",x"0FD03",x"0FCE3",x"0F4A3",x"0F463",x"0EC44",x"0EC67",x"0E52D",x"0DE55",
									 x"0E73B",x"0EF7D",x"0F7BE",x"0FFFF",x"10005",x"0FFFF",x"10006",x"0FFDF",x"0EF9D",x"0E73B",
									 x"0E678",x"0E570",x"0ECA9",x"0EC65",x"0F463",x"0F4A3",x"0F4C3",x"0FD03",x"0FD23",x"0FD64",
									 x"10000",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FDE5",x"10001",x"0FE05",x"10002",x"0FE25",
									 x"1000B",x"0FE45",x"10000",x"0FE46",x"10001",x"0FE26",x"0F606",x"0E565",x"0CCC4",x"0C4A4",
									 x"0C4C4",x"0CD04",x"0E585",x"0EDC6",x"0F605",x"0FE46",x"0FE65",x"0FE66",x"0FE85",x"10000",
									 x"0FE65",x"10023",x"0FE85",x"1002D",x"0FE65",x"1001A",x"0FE45",x"10000",x"0FE65",x"10002",
									 x"0FE45",x"0FE65",x"10000",x"0FE85",x"10004",x"0FE66",x"0FE46",x"0F627",x"0EDC6",x"0DD65",
									 x"0D504",x"0C4A4",x"10000",x"0CCE4",x"0DD65",x"0EDE6",x"0FE46",x"10001",x"0FE25",x"10010",
									 x"0FE05",x"10001",x"0FDE5",x"10001",x"0FDC5",x"0FDA5",x"0FDA4",x"0FD84",x"0FD64",x"10000",
									 x"0FD23",x"0FD03",x"0FCE3",x"0F4A3",x"0F463",x"0EC66",x"0EC89",x"0E54F",x"0DE76",x"0E73B",
									 x"0EF7D",x"0FFDF",x"0FFFF",x"10005",x"0FFFF",x"10006",x"0FFDF",x"0EF9E",x"0E73C",x"0E699",
									 x"0EDB2",x"0ECCA",x"0EC86",x"0F463",x"0F483",x"0F4A3",x"0FCE3",x"0FD23",x"0FD44",x"0FD64",
									 x"0FD84",x"10000",x"0FDA4",x"0FDC4",x"0FDC5",x"0FDE5",x"10000",x"0FE05",x"10002",x"0FE25",
									 x"1000B",x"0FE45",x"0FE46",x"10001",x"0FE26",x"0E584",x"0CCA5",x"0A382",x"08280",x"07A60",
									 x"08280",x"08AE1",x"0A382",x"0B402",x"0C4A3",x"0D524",x"0E584",x"0EDE5",x"0F645",x"0FE85",
									 x"10002",x"0FE65",x"10003",x"0FE85",x"0FE65",x"10019",x"0FE85",x"10033",x"0FE65",x"10019",
									 x"0FE85",x"10006",x"0FE65",x"0FE45",x"0F605",x"0E5A4",x"0D524",x"0CCC5",x"0B403",x"09B62",
									 x"092E2",x"08281",x"07A60",x"082A0",x"09B42",x"0C484",x"0EDE6",x"0FE26",x"0FE46",x"0FE25",
									 x"1000F",x"0FE05",x"10001",x"0FDE5",x"10002",x"0FDC5",x"0FDA5",x"0FDA4",x"0FD84",x"0FD64",
									 x"0FD43",x"0F523",x"0F503",x"0F4C3",x"0F483",x"0F464",x"0EC66",x"0ECAA",x"0E590",x"0E697",
									 x"0E73C",x"0F79E",x"0FFDF",x"0FFFF",x"10005",x"0FFFF",x"10006",x"0FFDF",x"0EF9E",x"0E73D",
									 x"0E6B9",x"0E5D3",x"0E4EC",x"0EC86",x"0F464",x"0F483",x"0F4A3",x"0FCE3",x"0FD23",x"0FD64",
									 x"10000",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"10000",x"0FDE5",x"10000",x"0FE05",x"10003",
									 x"0FE25",x"10008",x"0FE45",x"0FE25",x"10000",x"0FE46",x"10000",x"0FE65",x"0F605",x"0C483",
									 x"09302",x"069E1",x"05100",x"10001",x"06141",x"06981",x"071E1",x"08281",x"09B42",x"0ABE2",
									 x"0C463",x"0D523",x"0E5A4",x"0EDC4",x"0EE04",x"0F645",x"0FE65",x"10000",x"0FEA6",x"0FEA5",
									 x"0FEC5",x"0FEA5",x"0FE86",x"10000",x"0FEA5",x"0FE85",x"10000",x"0FE65",x"10004",x"0FE64",
									 x"0FE65",x"10008",x"0FE85",x"10039",x"0FE65",x"10003",x"0FE85",x"0FE65",x"0FE85",x"10001",
									 x"0FE66",x"0FE65",x"0FE85",x"0FE65",x"10006",x"0FE85",x"10000",x"0FEA5",x"10002",x"0FEA6",
									 x"10000",x"0FE86",x"0FE65",x"0FE25",x"0F605",x"0EDC4",x"0E584",x"0D524",x"0C4A3",x"0ABE2",
									 x"09B41",x"08281",x"07201",x"06180",x"05961",x"05121",x"05100",x"05101",x"06161",x"08AE2",
									 x"0CCE5",x"0E5C5",x"0FE65",x"0FE44",x"0FE45",x"0FE25",x"10002",x"0FE45",x"10001",x"0FE25",
									 x"10006",x"0FE05",x"10002",x"0FDE5",x"10000",x"0FDC5",x"0FDC4",x"0FDA5",x"0FDA4",x"0FD84",
									 x"0FD64",x"0F543",x"0F523",x"0F503",x"0F4C3",x"0F483",x"0F463",x"0F466",x"0E4CB",x"0E5B2",
									 x"0E6B8",x"0E71B",x"0F79E",x"0FFDF",x"0FFFF",x"10005",x"0FFFF",x"10006",x"0FFDF",x"0F79E",
									 x"0EF5D",x"0EEDA",x"0E614",x"0E50D",x"0EC87",x"0EC44",x"0F483",x"0F4A3",x"0F4E3",x"0FD23",
									 x"0FD44",x"0FD64",x"0FD84",x"0FDA4",x"10001",x"0FDC4",x"0FDE5",x"10001",x"0FE05",x"10002",
									 x"0FE25",x"1000B",x"0FE46",x"0FE65",x"0FE64",x"0E5A5",x"0A362",x"06180",x"048A0",x"03840",
									 x"04060",x"04080",x"04060",x"10001",x"050E0",x"06980",x"07A21",x"08AA2",x"0A364",x"0B404",
									 x"0C464",x"0CCC4",x"0DD64",x"0EDC4",x"0EE05",x"0F646",x"0F685",x"0FEA5",x"0FEC5",x"0FEA5",
									 x"0FEA6",x"10001",x"0FE86",x"0FEA6",x"10000",x"0FE85",x"10001",x"0FE84",x"0FE64",x"10000",
									 x"0FE65",x"0FE66",x"0FE65",x"10005",x"0FE85",x"10029",x"0FEA5",x"10001",x"0FE85",x"1000A",
									 x"0FE65",x"10007",x"0FE85",x"1000A",x"0FEA5",x"10002",x"0FEA6",x"10000",x"0FE85",x"0FE65",
									 x"0F665",x"0F625",x"0E5A5",x"0DD65",x"0D505",x"0C464",x"0ABC2",x"0A362",x"092E3",x"07A21",
									 x"06180",x"050E0",x"04060",x"03840",x"04080",x"04060",x"10000",x"03840",x"03820",x"061A0",
									 x"0AC03",x"0D544",x"0FE65",x"10000",x"0FE45",x"0FE25",x"1000D",x"0FE05",x"10002",x"0FDE5",
									 x"0FDE4",x"0FDC4",x"0FDA4",x"10000",x"0FD84",x"10000",x"0FD64",x"0F543",x"0F523",x"0F4E3",
									 x"0F4C3",x"0F482",x"0EC43",x"0EC87",x"0E4EC",x"0E5F3",x"0E6B9",x"0E73C",x"0F79E",x"0FFDF",
									 x"0FFFF",x"10005",x"0FFFF",x"10007",x"0F7BE",x"0EF5D",x"0E6FB",x"0E656",x"0E54E",x"0ECA9",
									 x"0EC44",x"0F463",x"0FCA3",x"0F4E3",x"0F503",x"0FD24",x"0FD44",x"0FD84",x"0FDA4",x"10001",
									 x"0FDC4",x"0FDE4",x"0FDE5",x"10000",x"0FE05",x"10002",x"0FE25",x"1000B",x"0FE45",x"0FE84",
									 x"0FE85",x"0D505",x"08261",x"050E0",x"04060",x"04881",x"050C1",x"050C0",x"10000",x"050C1",
									 x"050A0",x"050C0",x"058E1",x"05900",x"050E0",x"06100",x"06940",x"071A0",x"08260",x"09B21",
									 x"0ABA2",x"0B402",x"0C4A4",x"0CD24",x"0D564",x"0DDA4",x"0EE04",x"0F645",x"0FE65",x"0FEA6",
									 x"0FEC6",x"10002",x"0FEA6",x"10001",x"0FE86",x"0FE66",x"0FE65",x"0FE85",x"10007",x"0FE84",
									 x"10000",x"0FE85",x"10017",x"0FEA5",x"10004",x"0FE85",x"10004",x"0FEA5",x"10007",x"0FE85",
									 x"10010",x"0FE84",x"10000",x"0FEA4",x"0FE85",x"0FE86",x"10000",x"0FEA6",x"10001",x"0FEC6",
									 x"10002",x"0FEA6",x"0F665",x"0F645",x"0EE05",x"0E5A4",x"0DD44",x"0CCE4",x"0C4A3",x"0B422",
									 x"0A382",x"09301",x"08281",x"071E0",x"06140",x"06120",x"05900",x"058E0",x"050C0",x"050A0",
									 x"050C1",x"050C0",x"050E0",x"050C1",x"050E1",x"048A1",x"03820",x"05100",x"09322",x"0C4A3",
									 x"0FE46",x"0FE65",x"0FE45",x"0FE25",x"1000D",x"0FE05",x"10002",x"0FDE5",x"0FDE4",x"0FDC4",
									 x"0FDA4",x"10000",x"0FD84",x"10000",x"0FD64",x"0F543",x"0F503",x"0F4E3",x"0F4A3",x"0F482",
									 x"0EC64",x"0ECA8",x"0E50E",x"0E635",x"0E6FA",x"0EF5D",x"0F79E",x"0FFDF",x"0FFFF",x"10005",
									 x"0FFFF",x"10007",x"0F79E",x"0EF7D",x"0E73C",x"0E698",x"0DD70",x"0E4CA",x"0EC65",x"0F463",
									 x"0F4A3",x"0F4C3",x"0F503",x"0FD24",x"0FD44",x"0FD64",x"0FDA4",x"10001",x"0FDC4",x"0FDE4",
									 x"10000",x"0FDE5",x"0FE05",x"10001",x"0FE25",x"10008",x"0FE45",x"0FE25",x"10001",x"0FE45",
									 x"0FE84",x"0FE65",x"0CCE5",x"07A42",x"048A0",x"04880",x"058E1",x"06120",x"10000",x"06141",
									 x"10001",x"06101",x"05901",x"058E0",x"050C0",x"050A0",x"10000",x"058C0",x"06120",x"06981",
									 x"071C2",x"07A01",x"08AA2",x"09302",x"09B62",x"0ABE2",x"0BC84",x"0CD03",x"0D543",x"0DDA4",
									 x"0E5E4",x"0E624",x"0EE44",x"0EE64",x"0F684",x"10000",x"0FE84",x"0FEA4",x"10000",x"0FEA5",
									 x"0FEC5",x"10001",x"0FEA4",x"10000",x"0FEA5",x"10018",x"0FE85",x"10003",x"0FEA5",x"10004",
									 x"0FE85",x"1000A",x"0FEA5",x"10005",x"0FE85",x"10000",x"0FEA5",x"10001",x"0FE85",x"10002",
									 x"0FEA5",x"10001",x"0FEC5",x"10000",x"0FEC4",x"10002",x"0FEA4",x"0FEA5",x"10000",x"0F684",
									 x"10000",x"0F665",x"0EE45",x"0EE05",x"0E5C5",x"0DDA5",x"0D564",x"0CCE3",x"0BC82",x"0B403",
									 x"0A363",x"092C2",x"08282",x"08222",x"071C1",x"06980",x"06120",x"058E0",x"050A0",x"05080",
									 x"050A0",x"058E0",x"05900",x"06120",x"06140",x"10001",x"05921",x"05920",x"050E1",x"04061",
									 x"05120",x"082C1",x"0BC63",x"0F626",x"0FE65",x"0FE45",x"0FE25",x"1000D",x"0FE05",x"10002",
									 x"0FDE5",x"10000",x"0FDC4",x"0FDA4",x"0FD84",x"10000",x"0FD64",x"0FD44",x"0F523",x"0F503",
									 x"0F4E3",x"0F4A3",x"0F463",x"0EC44",x"0E4C9",x"0DD4F",x"0E656",x"0E71B",x"0EF7D",x"0F79E",
									 x"0FFFF",x"10006",x"0FFFF",x"10007",x"0F7BE",x"0EF7D",x"0E75D",x"0E6B9",x"0E5B2",x"0E4EB",
									 x"0EC45",x"0F463",x"0F483",x"0F4C3",x"0FD03",x"0FD24",x"0FD44",x"0FD84",x"0FDA4",x"10001",
									 x"0FDC4",x"0FDE4",x"10001",x"0FE04",x"0FE05",x"10000",x"0FE25",x"10005",x"0FE45",x"10006",
									 x"0FEA5",x"0FE85",x"0CCE5",x"07A41",x"04880",x"10000",x"06101",x"06120",x"06940",x"06960",
									 x"06940",x"06960",x"06940",x"10000",x"06941",x"06120",x"10001",x"05900",x"10000",x"058E1",
									 x"058C0",x"10000",x"058E0",x"05920",x"06160",x"071E0",x"08A82",x"09302",x"0A382",x"0ABE3",
									 x"0BC43",x"0C4A3",x"0D524",x"0DD64",x"0E5C4",x"0EE04",x"0F645",x"0F685",x"0FEA5",x"0FEC5",
									 x"0FEC6",x"10000",x"0FEE6",x"10001",x"0FEC6",x"10000",x"0FEC5",x"0FEA5",x"10002",x"0FEA4",
									 x"10000",x"0FEC4",x"10001",x"0FEC5",x"10000",x"0FEA4",x"10003",x"0FEA5",x"10001",x"0FEC5",
									 x"10000",x"0FEA5",x"10001",x"0FEA4",x"0FEA5",x"10013",x"0FEA4",x"10004",x"0FEA5",x"10001",
									 x"0FEA4",x"0FEA5",x"10004",x"0FEC5",x"10001",x"0FEE6",x"10003",x"0FEC6",x"0FEA5",x"0FE85",
									 x"0F645",x"0EE04",x"0E5C4",x"0DD64",x"0D505",x"0C484",x"0BC24",x"0B404",x"0A363",x"09302",
									 x"08281",x"07A01",x"06160",x"058E0",x"050A0",x"050C0",x"10000",x"058E0",x"10000",x"06100",
									 x"06101",x"06121",x"06940",x"10001",x"07160",x"10000",x"06960",x"06940",x"10000",x"06140",
									 x"05900",x"04880",x"05940",x"08AE2",x"0BC63",x"0F625",x"0FE65",x"0FE45",x"10000",x"0FE25",
									 x"10000",x"0FE45",x"0FE25",x"10009",x"0FE05",x"10002",x"0FDE5",x"0FDE4",x"0FDC4",x"0FDA4",
									 x"0FD84",x"10000",x"0FD64",x"0FD44",x"0FD24",x"0F503",x"0F4C3",x"0F483",x"0F462",x"0EC44",
									 x"0E4EA",x"0DD91",x"0DE78",x"0E73C",x"0EF7E",x"0F7BE",x"0FFFF",x"10006",x"0FFFF",x"10007",
									 x"0FFBE",x"0F79D",x"0E75D",x"0DEDA",x"0E5F4",x"0ED2D",x"0EC66",x"0F463",x"0F483",x"0F4A3",
									 x"0FCE3",x"0FD24",x"0FD44",x"0FD84",x"0FDA4",x"10001",x"0FDC4",x"0FDE4",x"10001",x"0FE04",
									 x"0FE05",x"10000",x"0FE25",x"10004",x"0FE45",x"10007",x"0FEA6",x"0FE86",x"0CD05",x"08261",
									 x"048A0",x"050A0",x"06921",x"07140",x"07160",x"07161",x"07160",x"10001",x"07181",x"10001",
									 x"06980",x"06960",x"06940",x"06140",x"06100",x"058E0",x"10000",x"050A0",x"10000",x"050C0",
									 x"05900",x"06120",x"06140",x"06160",x"06980",x"071C0",x"08240",x"08AA1",x"09B01",x"0A362",
									 x"0ABC3",x"0BC23",x"0C483",x"0CD04",x"0D544",x"0D583",x"0DDC4",x"0E604",x"0EE25",x"0EE45",
									 x"0F665",x"10000",x"0FE86",x"0FEA6",x"0FEC6",x"0FEE6",x"10000",x"0FF05",x"1000A",x"0FEE5",
									 x"10000",x"0FEC5",x"1001A",x"0FEE5",x"10004",x"0FF06",x"10004",x"0FEE6",x"0FEC5",x"10001",
									 x"0FEA5",x"0F685",x"0F665",x"0EE45",x"0EE25",x"0E605",x"0E5C4",x"0DDA4",x"0D544",x"0CCE4",
									 x"0C4A4",x"0BC43",x"0B403",x"0A362",x"09AE1",x"09280",x"08220",x"071A0",x"071A1",x"06141",
									 x"10000",x"06120",x"05900",x"050E1",x"050C0",x"10001",x"058E0",x"06100",x"06120",x"06940",
									 x"06960",x"07180",x"07161",x"07181",x"10000",x"07160",x"10001",x"07140",x"06941",x"06940",
									 x"06121",x"050A1",x"06140",x"08B02",x"0BC83",x"0F645",x"0FE65",x"0FE45",x"10000",x"0FE25",
									 x"0FE45",x"10000",x"0FE25",x"10009",x"0FE05",x"10001",x"0FDE5",x"10000",x"0FDC4",x"10000",
									 x"0FDA4",x"0FD84",x"10000",x"0FD64",x"0FD44",x"0FD24",x"0F503",x"0F4C3",x"0F483",x"0F462",
									 x"0EC65",x"0E52B",x"0DDD2",x"0DEB8",x"0E73C",x"0F79E",x"0F7BE",x"0FFFF",x"10006",x"0FFFF",
									 x"10007",x"0FFDF",x"0F79E",x"0EF7C",x"0E6DB",x"0DE16",x"0E54E",x"0EC87",x"0F443",x"0F483",
									 x"0F4A3",x"0FCE4",x"0FD24",x"0FD43",x"0FD64",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FDE4",
									 x"0FDE5",x"10000",x"0FE05",x"10000",x"0FE25",x"0FE05",x"0FE25",x"10002",x"0FE45",x"10007",
									 x"0FE66",x"0FEC6",x"0FEA6",x"0D565",x"08AC1",x"058E0",x"10000",x"06941",x"07140",x"07160",
									 x"10000",x"07980",x"10000",x"07981",x"10000",x"07980",x"10000",x"07180",x"07160",x"10001",
									 x"06960",x"06940",x"07161",x"06940",x"10000",x"06120",x"05900",x"050C0",x"050A0",x"10000",
									 x"04880",x"10000",x"048A0",x"050E0",x"05940",x"06180",x"071E0",x"07A21",x"08261",x"08AA1",
									 x"092E1",x"09B41",x"0A382",x"0ABE2",x"0B443",x"0C4A3",x"0CCE4",x"0D544",x"0DD85",x"0DDA4",
									 x"0E5E3",x"0E623",x"0EE64",x"10000",x"0EE84",x"0F6C5",x"0F6C4",x"0F6E5",x"10000",x"0FEC5",
									 x"0F6C5",x"0F6C4",x"0FEC5",x"10001",x"0FEE5",x"10002",x"0FEE6",x"0FEE5",x"0FEC5",x"10002",
									 x"0FEE5",x"0FEC5",x"10000",x"0FEE5",x"10004",x"0FEC4",x"0FEC5",x"10009",x"0F6C5",x"0FEC5",
									 x"10000",x"0F6C5",x"0F6C4",x"10000",x"0F6C5",x"0F6A4",x"0F6A5",x"0EE85",x"10000",x"0EE44",
									 x"0EE43",x"0E604",x"0DDC4",x"0DD84",x"0D544",x"0CD04",x"0C4A3",x"0BC63",x"0AC03",x"0A382",
									 x"09B42",x"09302",x"08AC1",x"08281",x"07A41",x"07201",x"069A0",x"05940",x"05100",x"048A0",
									 x"04880",x"10000",x"050A0",x"10000",x"058C0",x"05900",x"05920",x"06140",x"06160",x"06960",
									 x"10002",x"07160",x"07180",x"10001",x"07981",x"10001",x"079A1",x"079A0",x"07981",x"07961",
									 x"07160",x"06921",x"058A0",x"06160",x"09B42",x"0C4C3",x"0F686",x"0FE85",x"0FE65",x"0FE25",
									 x"10000",x"0FE45",x"10000",x"0FE25",x"10001",x"0FE24",x"0FE25",x"10004",x"0FE05",x"10001",
									 x"0FDE5",x"10001",x"0FDC4",x"0FDA4",x"10000",x"0FD84",x"10000",x"0FD64",x"0FD43",x"0FD23",
									 x"0FCE3",x"0F4A3",x"0F483",x"0F462",x"0EC66",x"0E54E",x"0D5F4",x"0DED9",x"0EF5D",x"0F79E",
									 x"0FFDF",x"0FFFF",x"10006",x"0FFFF",x"10007",x"0FFDF",x"0F79E",x"0EF7D",x"0DEDB",x"0DE37",
									 x"0ED90",x"0ECA8",x"0F444",x"0F483",x"0F4A3",x"0FCE4",x"0FD24",x"0FD43",x"0FD64",x"0FD84",
									 x"0FDA4",x"10000",x"0FDC4",x"0FDE5",x"10001",x"0FE05",x"10000",x"0FE25",x"10004",x"0FE45",
									 x"10007",x"0FE66",x"0FEC6",x"10000",x"0DD85",x"09321",x"06140",x"06100",x"06940",x"07161",
									 x"07981",x"079A1",x"079A0",x"10002",x"07180",x"10000",x"07160",x"10000",x"07180",x"10000",
									 x"06960",x"10000",x"07161",x"06960",x"10001",x"06140",x"06121",x"10000",x"06100",x"05900",
									 x"10005",x"05920",x"05940",x"10000",x"06161",x"06181",x"069A0",x"07200",x"08261",x"08AE1",
									 x"09321",x"09B62",x"0A3A2",x"0ABE3",x"0B443",x"0BC84",x"0BCA3",x"0C4C3",x"0C504",x"0CD44",
									 x"0D584",x"0D5A4",x"0DDC4",x"0DDC3",x"0E5E4",x"0E624",x"0EE44",x"0EE64",x"10000",x"0F684",
									 x"0F685",x"10000",x"0F6A5",x"0FEA5",x"0FEC5",x"10002",x"0FEE5",x"10000",x"0FF05",x"10005",
									 x"0FEE5",x"0FEC5",x"0FEE6",x"0FEC6",x"10000",x"0FEA5",x"0FE85",x"10001",x"0F685",x"0F664",
									 x"10001",x"0EE64",x"0E644",x"0E624",x"0E604",x"0DDC4",x"0DDA4",x"0D5A4",x"0D564",x"0CD44",
									 x"0C503",x"0C4E3",x"0BCA3",x"0BC83",x"0B443",x"0AC02",x"0A3A2",x"09B82",x"09321",x"08AC0",
									 x"08260",x"07A21",x"069C1",x"06161",x"06141",x"05920",x"10001",x"05921",x"05900",x"10001",
									 x"058E0",x"10000",x"05900",x"10000",x"06100",x"06120",x"06140",x"06960",x"10001",x"07180",
									 x"06981",x"06960",x"10000",x"07180",x"10001",x"07980",x"10001",x"079A1",x"10000",x"079A0",
									 x"07980",x"07981",x"07980",x"06921",x"058A0",x"06981",x"0A383",x"0CD24",x"0FEA6",x"0FE85",
									 x"0FE45",x"0FE25",x"10000",x"0FE45",x"10003",x"0FE25",x"10005",x"0FE05",x"10001",x"0FDE5",
									 x"10000",x"0FDC4",x"10001",x"0FDA4",x"0FD84",x"10000",x"0FD64",x"0FD43",x"0FD23",x"0FCE3",
									 x"0F4A3",x"0F483",x"0F463",x"0EC87",x"0E58F",x"0DE36",x"0DEDA",x"0EF5D",x"0F7BF",x"0FFDF",
									 x"0FFFF",x"10006",x"0FFFF",x"10007",x"0FFDF",x"0F7BE",x"0EF7D",x"0DEFB",x"0DE78",x"0E5D1",
									 x"0E4C9",x"0EC44",x"0F463",x"0FCA3",x"0FCC4",x"0FD04",x"0FD23",x"0FD64",x"0FD84",x"0FDA4",
									 x"10000",x"0FDC4",x"0FDE5",x"10001",x"0FE05",x"10000",x"0FE25",x"0FE05",x"0FE25",x"10002",
									 x"0FE45",x"10008",x"0FEC6",x"0FEC5",x"0E5C5",x"09B82",x"069A0",x"06140",x"06940",x"07981",
									 x"079A1",x"079A0",x"079C0",x"081C0",x"079C0",x"079A0",x"10001",x"071A0",x"07180",x"07160",
									 x"10000",x"06940",x"06961",x"10000",x"06981",x"06980",x"10000",x"06960",x"10003",x"06961",
									 x"06140",x"06120",x"05900",x"10000",x"058E0",x"050C0",x"10000",x"048A0",x"10001",x"050C0",
									 x"05100",x"05940",x"06160",x"06980",x"069A0",x"071C1",x"07201",x"07A22",x"07A42",x"08262",
									 x"08282",x"08AC2",x"09303",x"09342",x"09B82",x"09BA2",x"0A3C2",x"0ABE2",x"0B443",x"0BC83",
									 x"0BCA3",x"0C4C3",x"0C4E3",x"0CCE3",x"0CD03",x"10000",x"0D523",x"0D544",x"10000",x"0D564",
									 x"0DD84",x"0DDA4",x"10000",x"0DDC4",x"10000",x"0E5C4",x"10002",x"0DDC4",x"0DDA5",x"10002",
									 x"0D584",x"0D544",x"0D524",x"10001",x"0CD03",x"0CCE3",x"10000",x"0C4C3",x"0BC83",x"0B462",
									 x"0B423",x"0ABE3",x"0A3C3",x"0A3A3",x"09B83",x"09342",x"08B02",x"08AC2",x"082A1",x"08261",
									 x"08262",x"07A21",x"07201",x"071E0",x"069C0",x"069A0",x"06160",x"05940",x"05900",x"050C0",
									 x"048A0",x"04880",x"10000",x"050A0",x"050C0",x"05900",x"05901",x"06120",x"06140",x"06961",
									 x"10001",x"06980",x"06960",x"10003",x"07180",x"06960",x"06961",x"06960",x"10000",x"07160",
									 x"07180",x"07980",x"10002",x"079A0",x"079A1",x"079C0",x"079A0",x"07981",x"07980",x"07141",
									 x"058A0",x"069A1",x"0ABE3",x"0D544",x"0FEC6",x"0FE85",x"0FE45",x"10000",x"0FE25",x"0FE45",
									 x"10003",x"0FE25",x"10005",x"0FE05",x"10001",x"0FDE5",x"10000",x"0FDC4",x"10001",x"0FDA4",
									 x"0FD84",x"10000",x"0FD64",x"0FD43",x"0FD03",x"0FCE3",x"0F4A3",x"0F483",x"0EC64",x"0E4A8",
									 x"0E5B1",x"0DE77",x"0DEFA",x"0EF5D",x"0F7BF",x"0FFDF",x"0FFFF",x"10006",x"0FFFF",x"10008",
									 x"0FFDF",x"0F79D",x"0E71C",x"0E6DA",x"0E634",x"0E4EB",x"0EC65",x"0EC63",x"0F4A3",x"0FCC4",
									 x"0FD03",x"0F523",x"0FD43",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"10000",x"0FDE5",x"10000",
									 x"0FE05",x"10000",x"0FE25",x"10004",x"0FE45",x"10005",x"0FE25",x"0FE24",x"0FE45",x"0FEA5",
									 x"0FEC5",x"0E605",x"0AC02",x"07A41",x"06960",x"06920",x"07161",x"079A1",x"081C1",x"081C0",
									 x"081A0",x"07980",x"079A0",x"079C2",x"07A02",x"079E3",x"079C2",x"07182",x"06961",x"06121",
									 x"10000",x"05920",x"05940",x"10000",x"06160",x"06980",x"10000",x"06960",x"10000",x"06981",
									 x"10000",x"06960",x"10000",x"06940",x"06140",x"10000",x"06160",x"10000",x"06140",x"10000",
									 x"05940",x"05920",x"10000",x"05900",x"10001",x"058E0",x"050E0",x"050C0",x"10001",x"048A0",
									 x"10000",x"050C0",x"05100",x"05920",x"05940",x"06140",x"06160",x"06180",x"069C0",x"07200",
									 x"07A41",x"07A40",x"10000",x"08260",x"10000",x"08280",x"10000",x"082A1",x"082C1",x"08AE1",
									 x"10000",x"09301",x"10000",x"09321",x"10007",x"09301",x"08AE1",x"08AC0",x"082C0",x"08281",
									 x"10000",x"08261",x"10000",x"08260",x"08240",x"07A60",x"07A40",x"07200",x"069E1",x"069A1",
									 x"06160",x"06140",x"05940",x"05900",x"050E0",x"10000",x"050C0",x"10002",x"050E0",x"10002",
									 x"05900",x"05920",x"10000",x"05940",x"06140",x"10000",x"06141",x"06140",x"06160",x"10002",
									 x"06961",x"10000",x"06960",x"10001",x"06160",x"10000",x"06960",x"10000",x"06940",x"06140",
									 x"10001",x"06120",x"06940",x"07181",x"079E2",x"07A02",x"07A03",x"079C2",x"07180",x"079A1",
									 x"079A0",x"081E0",x"081C0",x"079A1",x"079A0",x"07161",x"058E0",x"07201",x"0B443",x"0DDA4",
									 x"0FEC6",x"0FE85",x"0FE45",x"10000",x"0FE25",x"0FE45",x"10006",x"0FE25",x"10002",x"0FE05",
									 x"10001",x"0FDE5",x"10000",x"0FDC4",x"10000",x"0FDA4",x"10000",x"0FD84",x"0FD64",x"0F564",
									 x"0F544",x"0FD03",x"0FCC3",x"0F4A3",x"0F463",x"0EC64",x"0E4AA",x"0EDF3",x"0E6B9",x"0DF1B",
									 x"0EF7D",x"0FFDF",x"10000",x"0FFFF",x"10006",x"0FFFF",x"10007",x"0FFDF",x"10000",x"0F79D",
									 x"0E73D",x"0E6FB",x"0E655",x"0E52C",x"0E466",x"0EC63",x"0F483",x"0FCC3",x"0FCE3",x"0F523",
									 x"0FD43",x"0FD64",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FDE4",x"0FDE5",x"0FE05",x"10001",
									 x"0FE25",x"10002",x"0FE45",x"10006",x"0FE44",x"0FE24",x"0FE45",x"0FE85",x"0FEC5",x"0EE45",
									 x"0B443",x"08AA1",x"071A0",x"06920",x"07961",x"07981",x"079A0",x"081A0",x"079A1",x"081E2",
									 x"08265",x"08AE7",x"08B29",x"0932A",x"08B09",x"082C8",x"07AA7",x"07266",x"07246",x"06A24",
									 x"061E3",x"061C1",x"06180",x"10000",x"06140",x"05920",x"10001",x"06140",x"10000",x"06160",
									 x"10000",x"06960",x"06980",x"10001",x"06981",x"06980",x"10000",x"06960",x"06160",x"06140",
									 x"06120",x"05920",x"10000",x"05900",x"10000",x"058E0",x"050E0",x"10000",x"050C0",x"10002",
									 x"058E0",x"10001",x"05900",x"05920",x"05940",x"06140",x"10001",x"06160",x"10002",x"06161",
									 x"10001",x"06181",x"069A1",x"1000B",x"06181",x"10000",x"06161",x"10005",x"06140",x"05920",
									 x"05900",x"10000",x"058E0",x"10000",x"050E0",x"050C0",x"10003",x"050E0",x"058E0",x"05900",
									 x"10000",x"05920",x"06120",x"06140",x"10000",x"06160",x"06960",x"06980",x"10003",x"06960",
									 x"10001",x"06161",x"06140",x"10000",x"05920",x"10000",x"05940",x"06140",x"06160",x"06981",
									 x"069A2",x"069C2",x"06A03",x"07225",x"07A66",x"07AA7",x"082C7",x"08B29",x"0936A",x"10000",
									 x"08AE8",x"08265",x"081E2",x"07980",x"079C0",x"10000",x"079A1",x"079A0",x"07160",x"06100",
									 x"07A21",x"0BC83",x"0E5C4",x"0FEC6",x"0FE85",x"0FE45",x"10000",x"0FE25",x"0FE45",x"10006",
									 x"0FE25",x"10002",x"0FE05",x"10001",x"0FDE5",x"10000",x"0FDC4",x"10000",x"0FDA4",x"10000",
									 x"0FD84",x"0FD64",x"0F564",x"0F544",x"0FCE3",x"0FCC3",x"0F483",x"0EC63",x"0EC85",x"0E4EC",
									 x"0EE55",x"0E6FB",x"0E73C",x"0F79D",x"0FFDE",x"0FFDF",x"0FFFF",x"10006",x"0FFFF",x"10008",
									 x"0FFDF",x"0F7BE",x"0E73D",x"0E71C",x"0E676",x"0E56E",x"0EC87",x"0EC64",x"0F462",x"0FCA3",
									 x"0FCE3",x"0F523",x"0FD43",x"0FD64",x"0FD84",x"10000",x"0FDA4",x"0FDC4",x"10000",x"0FDE4",
									 x"0FDE5",x"0FE05",x"10000",x"0FE25",x"10002",x"0FE45",x"10001",x"0FE44",x"0FE45",x"0FE65",
									 x"0FE44",x"10001",x"0FE24",x"0FE45",x"0FE85",x"0FEC5",x"0F666",x"0BCA3",x"09302",x"071E0",
									 x"06120",x"07161",x"081C1",x"081E0",x"079A0",x"071A1",x"08265",x"0936A",x"0A44E",x"0A490",
									 x"0ACB1",x"0A490",x"0A46F",x"09C4E",x"08BED",x"083AB",x"08349",x"07AC6",x"07265",x"06A03",
									 x"069C2",x"06182",x"05962",x"05942",x"05940",x"10000",x"06160",x"10001",x"06140",x"10001",
									 x"06941",x"10001",x"06961",x"10001",x"06960",x"10000",x"06160",x"10001",x"06980",x"06180",
									 x"06160",x"10001",x"06140",x"10001",x"06141",x"06120",x"06140",x"10000",x"05940",x"05920",
									 x"10003",x"05900",x"10001",x"05100",x"10000",x"050E0",x"10010",x"05100",x"10003",x"05920",
									 x"10001",x"05900",x"05920",x"10000",x"06120",x"06141",x"10001",x"06140",x"10000",x"06160",
									 x"10002",x"06180",x"06160",x"10000",x"06960",x"10001",x"06940",x"06961",x"06960",x"10000",
									 x"06160",x"06140",x"10002",x"06141",x"06140",x"06160",x"05941",x"10000",x"05962",x"06182",
									 x"061A2",x"069E3",x"07265",x"07AC6",x"08328",x"08B8C",x"093CD",x"0940E",x"09C4F",x"0A4B1",
									 x"10001",x"09C0E",x"09349",x"08A64",x"079A0",x"081C0",x"079A0",x"079A1",x"079A0",x"07160",
									 x"06120",x"08A81",x"0CCE4",x"0E5E4",x"0FEC5",x"0FE85",x"0FE45",x"10000",x"0FE25",x"0FE45",
									 x"10006",x"0FE25",x"10002",x"0FE05",x"10001",x"0FDE5",x"10000",x"0FDC4",x"10000",x"0FDA4",
									 x"10000",x"0FD84",x"0FD64",x"0F544",x"0F523",x"0FCE3",x"0FCA3",x"0F463",x"0EC63",x"0ECA6",
									 x"0E52D",x"0EE56",x"0E6FB",x"0E75D",x"0F79D",x"0FFDE",x"0FFFF",x"10007",x"0FFFF",x"10008",
									 x"0FFDE",x"0F7BF",x"0EF5E",x"0E71B",x"0E6B8",x"0DDB1",x"0E4A9",x"0F444",x"0FC42",x"0FCA2",
									 x"0F4E3",x"0F503",x"0FD23",x"0FD64",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"10000",x"0FDE5",
									 x"10000",x"0FE05",x"10001",x"0FE25",x"10001",x"0FE45",x"10004",x"0FE65",x"0FE45",x"10002",
									 x"0FE65",x"0FEA5",x"0FEA6",x"0CD24",x"0A382",x"079E1",x"06100",x"07180",x"079C0",x"10000",
									 x"071A0",x"071C2",x"08B09",x"0A491",x"0B595",x"0B5D7",x"0BDD7",x"10000",x"0BDB6",x"0BDD6",
									 x"0B5B5",x"0AD74",x"0AD12",x"0ACAF",x"0A44E",x"09C0D",x"093AC",x"0934B",x"08B2A",x"0832A",
									 x"07AE8",x"07A85",x"07243",x"07201",x"069C1",x"06181",x"06140",x"05920",x"05900",x"058E0",
									 x"05901",x"05900",x"05920",x"05900",x"05920",x"06140",x"10000",x"06160",x"06180",x"10000",
									 x"061A0",x"10000",x"061C0",x"061A0",x"06980",x"10000",x"06960",x"06180",x"10003",x"06160",
									 x"05960",x"05940",x"10000",x"06140",x"10005",x"05940",x"06140",x"05940",x"10003",x"05920",
									 x"05940",x"10001",x"06140",x"05940",x"10000",x"06140",x"10007",x"06160",x"10002",x"06180",
									 x"06961",x"10000",x"06981",x"10000",x"06980",x"10000",x"069A0",x"06180",x"10000",x"06160",
									 x"10001",x"06140",x"10000",x"05920",x"06140",x"05920",x"05900",x"10002",x"05920",x"05940",
									 x"069A1",x"069C1",x"06A02",x"07243",x"072A6",x"07AE8",x"0832A",x"0836A",x"08B6B",x"08B8B",
									 x"09BED",x"0A46F",x"0A4B0",x"0AD32",x"0B575",x"0BDB6",x"10000",x"0B5B6",x"10000",x"0B5D7",
									 x"10000",x"0B554",x"0A46F",x"08B08",x"079C1",x"079C0",x"071A0",x"079C1",x"07961",x"07141",
									 x"07180",x"09B22",x"0D564",x"0EE44",x"0FEC5",x"0FE85",x"0FE45",x"0FE25",x"0FE45",x"10007",
									 x"0FE25",x"10002",x"0FE05",x"10001",x"0FDE5",x"10000",x"0FDE4",x"0FDC4",x"0FDA4",x"10000",
									 x"0FD84",x"0FD64",x"0FD44",x"0F523",x"0F503",x"0F4A3",x"0F463",x"0F444",x"0ECA8",x"0E570",
									 x"0E678",x"0DF1B",x"0E77E",x"0F7BE",x"0FFFE",x"0FFFF",x"10007",x"0FFFF",x"10008",x"0FFDE",
									 x"0F7DF",x"0EF7E",x"0E71B",x"0E6B8",x"0E5F3",x"0E4CB",x"0EC65",x"0F442",x"0F482",x"0F4C3",
									 x"0F503",x"0FD23",x"0FD44",x"0FD84",x"10000",x"0FDA4",x"0FDC4",x"10000",x"0FDE5",x"10000",
									 x"0FE05",x"10001",x"0FE25",x"10004",x"0FE45",x"10001",x"0FE65",x"0FE45",x"0FE65",x"0FE45",
									 x"10000",x"0FE65",x"0FE85",x"0FEC6",x"0D584",x"0AC03",x"07A21",x"060E0",x"07181",x"079C0",
									 x"10000",x"07180",x"071C3",x"0936B",x"0B533",x"0BE18",x"10000",x"0BDF9",x"0BE19",x"0C639",
									 x"10000",x"0C638",x"0BE18",x"0C5F7",x"0BDB5",x"0BD94",x"0B553",x"0B533",x"0AD13",x"0ACF3",
									 x"0ACD1",x"0A46F",x"09C0D",x"093AB",x"08B48",x"082E7",x"07A85",x"07245",x"06A24",x"06A04",
									 x"061E4",x"061C4",x"061A3",x"069A2",x"06182",x"06981",x"06180",x"06160",x"10001",x"06140",
									 x"10001",x"06160",x"05940",x"06140",x"10001",x"06160",x"10002",x"06140",x"06160",x"10009",
									 x"06180",x"06181",x"10001",x"06180",x"10000",x"061A0",x"06180",x"10002",x"06181",x"10000",
									 x"06160",x"10002",x"06961",x"10002",x"06960",x"06141",x"10000",x"06140",x"06141",x"10000",
									 x"06140",x"10009",x"06160",x"10001",x"06180",x"061A0",x"061A1",x"061C2",x"061C3",x"10000",
									 x"069E4",x"06A05",x"10000",x"07245",x"07AA6",x"07AE6",x"08328",x"08BAA",x"09C2D",x"0A490",
									 x"0A4D2",x"0ACF3",x"0AD13",x"0AD33",x"0B554",x"0B595",x"0BDD5",x"0BDF6",x"0C617",x"0C638",
									 x"10000",x"0C618",x"0BE18",x"10000",x"0BE39",x"0BDD6",x"0ACF1",x"09389",x"07A01",x"079C0",
									 x"071A0",x"079C0",x"07140",x"07141",x"079E1",x"0A3A3",x"0DDC5",x"0F665",x"0FEA4",x"0FE64",
									 x"0FE45",x"10009",x"0FE25",x"10002",x"0FE05",x"10000",x"0FDE5",x"10000",x"0FDE4",x"0FDC4",
									 x"10000",x"0FDA4",x"0FD84",x"0FD64",x"0FD44",x"0FD23",x"0F503",x"0F4E2",x"0F4A3",x"0F464",
									 x"0EC45",x"0ECC9",x"0E5B2",x"0E698",x"0E71B",x"0EF7E",x"0F7DF",x"0FFFE",x"0FFFF",x"10007",
									 x"0FFFF",x"10009",x"0F7DF",x"0EF7E",x"0E71C",x"0DEB9",x"0E635",x"0E50D",x"0EC67",x"0F443",
									 x"0F483",x"0F4C3",x"0FD03",x"0FD23",x"0FD44",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"10000",
									 x"0FDE5",x"10000",x"0FE05",x"10001",x"0FE25",x"10004",x"0FE45",x"10001",x"0FE65",x"0FE45",
									 x"10002",x"0FE65",x"0FEA5",x"0FEC6",x"0DDC4",x"0B463",x"07A40",x"058E0",x"07181",x"079C0",
									 x"071C0",x"07161",x"069C3",x"0938C",x"0B554",x"0BE38",x"0B618",x"0B5F8",x"0BDF8",x"0BE19",
									 x"0BE18",x"10001",x"0C618",x"10000",x"0C638",x"0BE18",x"10000",x"0C638",x"10000",x"0C617",
									 x"0BDD6",x"0BD95",x"0B553",x"0ACF1",x"0ACB0",x"0A46F",x"09C4F",x"09C0E",x"0940D",x"093ED",
									 x"093AC",x"08B6A",x"08B49",x"08307",x"07AA5",x"07263",x"07222",x"069E2",x"06181",x"06161",
									 x"06141",x"05921",x"05920",x"10000",x"05100",x"10000",x"05120",x"10001",x"05920",x"10001",
									 x"05940",x"10000",x"06140",x"10001",x"06160",x"10008",x"06180",x"10004",x"06160",x"10004",
									 x"06140",x"10007",x"06120",x"05920",x"05900",x"10000",x"05100",x"05900",x"05100",x"10000",
									 x"05120",x"05920",x"05940",x"05941",x"06161",x"06181",x"069C1",x"06A02",x"07243",x"07284",
									 x"07AE6",x"08349",x"0838B",x"08BAC",x"093CD",x"09BEE",x"09C0E",x"09C2E",x"0A46F",x"0A4AF",
									 x"0A4D0",x"0AD32",x"0BD94",x"0BDB6",x"0BDF8",x"10000",x"0C618",x"0C638",x"0C618",x"0C617",
									 x"10001",x"0C618",x"10000",x"0BE18",x"10000",x"0BDF8",x"0B5F8",x"0B618",x"0B5B6",x"0ACF1",
									 x"0938A",x"071E2",x"071A0",x"10000",x"079C0",x"06940",x"06941",x"07A20",x"0AC22",x"0E625",
									 x"0F685",x"0FE84",x"0FE65",x"0FE45",x"10009",x"0FE25",x"10002",x"0FE05",x"10000",x"0FDE5",
									 x"0FDE4",x"0FDC4",x"10001",x"0FDA4",x"0FD84",x"0FD64",x"0FD43",x"0FD23",x"0F503",x"0F4E3",
									 x"0F4A3",x"0F444",x"0EC66",x"0E4EB",x"0E5F4",x"0DE99",x"0E71B",x"0EF7E",x"0F7DF",x"0FFFE",
									 x"0FFFF",x"10007",x"0FFFF",x"10009",x"0F7DF",x"0EF9E",x"0E73C",x"0DEDA",x"0E678",x"0DD70",
									 x"0E4A9",x"0EC44",x"0F483",x"0F4C3",x"0F4E2",x"0F503",x"0FD44",x"0FD64",x"0FD84",x"0FDA4",
									 x"0FDC4",x"10000",x"0FDE4",x"0FDE5",x"10000",x"0FE05",x"10000",x"0FE25",x"10004",x"0FE45",
									 x"10006",x"0FE65",x"0FE84",x"0FEE6",x"0E624",x"0C4E3",x"082A1",x"05900",x"06961",x"071C1",
									 x"10000",x"06960",x"069C3",x"08B6B",x"0AD33",x"0BE17",x"0BE18",x"0BDF7",x"10000",x"0BE18",
									 x"0BE17",x"0BE18",x"0C638",x"10000",x"0C639",x"0CE3A",x"0CE5A",x"10000",x"0CE7A",x"0CE9A",
									 x"0CE7A",x"10000",x"0CE79",x"0C638",x"0C617",x"0C5F7",x"0C5F8",x"0C5D7",x"10000",x"0C5B6",
									 x"0BDB6",x"0B594",x"0AD52",x"0AD11",x"0A4CF",x"09C6C",x"0940A",x"093EA",x"0938A",x"08B29",
									 x"08309",x"082C9",x"082A8",x"07AA8",x"10000",x"07287",x"10000",x"06A66",x"10000",x"06A45",
									 x"06A24",x"10000",x"06A23",x"06A02",x"061E1",x"061C0",x"069A0",x"061A0",x"069A0",x"10001",
									 x"061A0",x"069A0",x"10000",x"06180",x"10000",x"06160",x"10000",x"06140",x"10000",x"05920",
									 x"05940",x"06140",x"06160",x"10000",x"06180",x"10001",x"061A0",x"10001",x"061C0",x"10003",
									 x"061C1",x"069C1",x"069E2",x"069E3",x"07224",x"10000",x"07245",x"06A46",x"07266",x"07287",
									 x"10000",x"07AA8",x"07AC8",x"10000",x"082C8",x"082E8",x"08B29",x"0936A",x"093AB",x"093EC",
									 x"09C2D",x"0A48F",x"0ACF2",x"0AD34",x"0B555",x"0BD95",x"0BDB6",x"0BDD6",x"0C5D6",x"0C5F7",
									 x"10000",x"0C617",x"0C637",x"0C638",x"0CE5A",x"0CE7A",x"0CE5A",x"0CE59",x"10001",x"0C638",
									 x"10001",x"0BE38",x"0BE18",x"0BDF8",x"10000",x"0BDD8",x"0BDF8",x"0BE38",x"0B5D6",x"0A4D1",
									 x"08B6A",x"061A1",x"069A0",x"069C0",x"071C1",x"06120",x"06961",x"08260",x"0BCC3",x"0F6A5",
									 x"0FEC5",x"0FE84",x"0FE45",x"10000",x"0FE44",x"0FE45",x"10007",x"0FE25",x"10002",x"0FE05",
									 x"10000",x"0FDE5",x"10000",x"0FDC4",x"10000",x"0FDA4",x"10000",x"0FD84",x"0FD64",x"0FD43",
									 x"0FD23",x"0F503",x"0F4E2",x"0F4A3",x"0EC65",x"0E487",x"0E54D",x"0E657",x"0E6DB",x"0E73B",
									 x"0F79E",x"0FFDF",x"0FFFE",x"0FFFF",x"10007",x"0FFFF",x"1000A",x"0F7BE",x"0E75D",x"0DEFC",
									 x"0E6BA",x"0DDB3",x"0E4CA",x"0EC45",x"0F483",x"0F4A2",x"0F4C2",x"0FD03",x"0FD24",x"0FD64",
									 x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FDE4",x"0FDE5",x"10000",x"0FE05",x"10000",x"0FE25",
									 x"10004",x"0FE45",x"10006",x"0FE44",x"0FE84",x"0FEE5",x"0EE64",x"0D584",x"09B62",x"06960",
									 x"06961",x"06980",x"071A1",x"06160",x"06181",x"07AE8",x"09CB0",x"0B5B5",x"0BDF7",x"0BE17",
									 x"0C617",x"10000",x"0C618",x"0C638",x"10001",x"0CE38",x"0CE59",x"10000",x"0CE39",x"0CE59",
									 x"10000",x"0CE7A",x"10000",x"0CE9A",x"10001",x"0D69B",x"10000",x"0D6BB",x"10000",x"0D6DB",
									 x"10000",x"0D6DA",x"0CEB9",x"0CE99",x"0CE78",x"0C636",x"0C616",x"0C615",x"0CDF5",x"0C5D5",
									 x"0C5B5",x"0C595",x"10000",x"0BD74",x"10001",x"0B554",x"0AD32",x"0AD11",x"0ACD0",x"0ACAF",
									 x"0A46E",x"09C2D",x"09C0B",x"093CA",x"093A9",x"09369",x"08B68",x"10001",x"08B48",x"10000",
									 x"08B28",x"08B27",x"08B07",x"08307",x"082E6",x"082C6",x"082A7",x"07A86",x"10002",x"07AA7",
									 x"082C6",x"082E7",x"08307",x"08B28",x"08B48",x"10000",x"08B68",x"10000",x"08368",x"08B68",
									 x"08B88",x"10000",x"08B89",x"093CA",x"09BEB",x"09C2C",x"0A46E",x"0ACAF",x"0ACD0",x"0ACF1",
									 x"0B512",x"0B533",x"0BD54",x"0BD75",x"0BD95",x"0BD94",x"10000",x"0BD95",x"0C5B5",x"0C5D6",
									 x"0CDF6",x"0CE17",x"0CE37",x"0CE58",x"0D679",x"0D67A",x"0D69B",x"0D6BA",x"10000",x"0D6DA",
									 x"0D6BA",x"0D69A",x"0CE9A",x"10000",x"0CE7A",x"10001",x"0CE59",x"0CE39",x"0CE38",x"0C638",
									 x"10001",x"0C618",x"0CE38",x"0C658",x"0C618",x"10000",x"0C5F8",x"10000",x"0BE18",x"0BE39",
									 x"0B5B6",x"09C90",x"07AE8",x"05960",x"069A0",x"069C0",x"071C1",x"06120",x"06960",x"08AE1",
									 x"0CD64",x"0F6E5",x"0FEE5",x"0FE84",x"0FE45",x"10000",x"0FE64",x"0FE45",x"10007",x"0FE25",
									 x"10002",x"0FE05",x"10000",x"0FDE5",x"10000",x"0FDC4",x"10000",x"0FDA4",x"10000",x"0FD84",
									 x"0FD44",x"0FD23",x"0FD03",x"0F4E2",x"0F4C2",x"0F483",x"0EC66",x"0E4A9",x"0E590",x"0E699",
									 x"0E6FC",x"0E73C",x"0F79E",x"0FFDF",x"0FFFF",x"10008",x"0FFFF",x"1000A",x"0F7DE",x"0EF7D",
									 x"0E71D",x"0E6FB",x"0DDF4",x"0E50C",x"0E465",x"0EC63",x"0F482",x"0FCC2",x"0F503",x"0FD23",
									 x"0FD44",x"0FD64",x"0FDA4",x"10000",x"0FDC4",x"0FDE5",x"10001",x"0FE05",x"10000",x"0FE25",
									 x"10004",x"0FE45",x"10007",x"0FE84",x"0FEC5",x"0EEA4",x"0DDE5",x"0A3E3",x"071E1",x"06961",
									 x"06960",x"069A1",x"06160",x"059A1",x"06A65",x"08C0D",x"0B553",x"0BDD6",x"0C618",x"10002",
									 x"0CE39",x"10000",x"0C638",x"0C658",x"0CE58",x"0CE59",x"0CE58",x"0CE78",x"0CE79",x"0CE7A",
									 x"10001",x"0CE9A",x"10001",x"0D6BA",x"0D6DA",x"0D6BA",x"10000",x"0D6BB",x"10000",x"0D6BA",
									 x"0D6BB",x"10003",x"0DEBA",x"0DEDB",x"0D6DB",x"10000",x"0D6FB",x"0DEFB",x"0DEDA",x"0D6DA",
									 x"10000",x"0D6B9",x"0D699",x"0D698",x"0D678",x"0CE37",x"0CE16",x"0CDD5",x"0CDD4",x"10000",
									 x"0C5B3",x"10001",x"0BDB3",x"10000",x"0BD93",x"0C593",x"10001",x"0C572",x"0BD72",x"0BD52",
									 x"0BD32",x"10003",x"0BD52",x"0BD72",x"0BD73",x"0C573",x"0C593",x"0C5B3",x"10002",x"0C593",
									 x"10000",x"0C5B3",x"10000",x"0C5D3",x"0C5D4",x"0CDF5",x"0CE16",x"0CE37",x"0D678",x"0D698",
									 x"0D699",x"0D6B9",x"0D6DA",x"0DEDB",x"0DEDC",x"0DEDB",x"0D6DB",x"10004",x"0D6BA",x"10002",
									 x"0D6BB",x"0DEDB",x"0D6BA",x"0D69A",x"0CEBA",x"0CE9A",x"10000",x"0CE7B",x"0D67B",x"0D69A",
									 x"10000",x"0D679",x"0CE58",x"10000",x"0CE59",x"10000",x"0C659",x"10000",x"0C639",x"10000",
									 x"0C658",x"0C638",x"10000",x"0C618",x"0C5F7",x"0C618",x"0BE39",x"0B575",x"0942F",x"07286",
									 x"05100",x"06160",x"069C0",x"069C1",x"06120",x"06980",x"09342",x"0D5E4",x"0FF25",x"0FEE5",
									 x"0FE64",x"0FE25",x"0FE45",x"0FE64",x"0FE45",x"10001",x"0FE65",x"0FE45",x"10003",x"0FE25",
									 x"10002",x"0FE05",x"10000",x"0FDE5",x"10000",x"0FDC4",x"10000",x"0FDA4",x"10000",x"0FD64",
									 x"0FD44",x"0FD23",x"0FD03",x"0F4C2",x"0F4A2",x"0EC63",x"0EC66",x"0E4EA",x"0E5D2",x"0E6DA",
									 x"0E71D",x"0EF7C",x"0FFBF",x"0FFFF",x"10009",x"0FFFF",x"1000A",x"0FFDF",x"0F79E",x"0E75D",
									 x"0E6FA",x"0DE15",x"0DD2E",x"0EC87",x"0F422",x"0F483",x"0F4C3",x"0F4E3",x"0FD03",x"0FD44",
									 x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"10000",x"0FDE4",x"0FE05",x"10001",x"0FE25",x"10001",
									 x"0FE45",x"10007",x"0FE44",x"0FE45",x"10000",x"0FE65",x"0FEA5",x"0F6A5",x"0EE65",x"0B483",
									 x"07A40",x"06940",x"06960",x"069A0",x"061A0",x"05980",x"059E3",x"0838A",x"0AD12",x"0BDD6",
									 x"0C639",x"10000",x"0C638",x"10000",x"0CE58",x"0CE38",x"0CE59",x"10002",x"0CE79",x"10002",
									 x"0D69A",x"10005",x"0D6BA",x"10002",x"0DEDA",x"0DEDB",x"10000",x"0DEFB",x"10001",x"0E71C",
									 x"10001",x"0E73C",x"10001",x"0EF3D",x"0E73D",x"0E73C",x"10000",x"0E71C",x"10001",x"0DEFB",
									 x"0DEDB",x"10000",x"0DEDA",x"0DEBA",x"10000",x"0D6BA",x"10004",x"0DEBA",x"0D6BA",x"10000",
									 x"0D6B9",x"10000",x"0D699",x"0D6B9",x"0D699",x"10004",x"0DE99",x"0DEBA",x"10004",x"0D6BA",
									 x"10000",x"0DEBA",x"10000",x"0DEDB",x"10001",x"0DEFB",x"10000",x"0DF1B",x"0E71C",x"0E73C",
									 x"10006",x"0E71C",x"0DF1C",x"0DEFC",x"0DEFB",x"10001",x"0DEDB",x"10000",x"0D6BB",x"0D6BA",
									 x"0D69A",x"10006",x"0D679",x"0CE79",x"10002",x"0CE59",x"10003",x"0C638",x"10001",x"0C617",
									 x"0C638",x"0BE18",x"0AD12",x"093AB",x"06A25",x"04920",x"06160",x"069C0",x"069A0",x"06160",
									 x"071E0",x"0A3C1",x"0E624",x"0FF25",x"0FEE5",x"0FE44",x"0FE45",x"10000",x"0FE65",x"10000",
									 x"0FE45",x"10000",x"0FE65",x"0FE45",x"10003",x"0FE25",x"10002",x"0FE05",x"10000",x"0FDE5",
									 x"0FDE4",x"0FDC4",x"0FDA4",x"10000",x"0FD83",x"0FD63",x"0FD43",x"0FD03",x"0FCE3",x"0F4A3",
									 x"0F482",x"0EC63",x"0E486",x"0E52D",x"0DDF4",x"0E6DA",x"0EF3C",x"0EF7D",x"0F7BF",x"0FFFF",
									 x"10009",x"0FFFF",x"1000A",x"0FFDF",x"0F79E",x"0EF5D",x"0E6FB",x"0DE36",x"0DD91",x"0ECC9",
									 x"0F443",x"0F463",x"0F4A3",x"0F4E3",x"0FD03",x"0FD23",x"0FD63",x"0FD84",x"0FDA4",x"10000",
									 x"0FDC4",x"0FDE4",x"0FE05",x"10001",x"0FE25",x"10001",x"0FE45",x"10007",x"0FE44",x"0FE45",
									 x"10000",x"0FE65",x"0FE85",x"0FEE5",x"0F6E6",x"0C544",x"082C2",x"06960",x"06140",x"061A0",
									 x"10000",x"05180",x"04981",x"06AC7",x"09CB0",x"0BDB6",x"0C639",x"10000",x"0C618",x"0C638",
									 x"0CE58",x"0C638",x"0CE59",x"10001",x"0CE79",x"10001",x"0D69A",x"10003",x"0D6BA",x"10001",
									 x"0DEDB",x"10004",x"0DEFB",x"10002",x"0E71C",x"10004",x"0E73C",x"10001",x"0E71C",x"0E73C",
									 x"0E73D",x"0EF5D",x"10007",x"0EF7D",x"10002",x"0F79D",x"1000B",x"0F77D",x"0F79D",x"10002",
									 x"0F77D",x"10000",x"0EF7D",x"10001",x"0EF5D",x"0EF7D",x"10000",x"0EF5D",x"10003",x"0E75C",
									 x"0E73C",x"10005",x"0E71C",x"0DF1C",x"0DF1B",x"0E71C",x"0DEFB",x"10001",x"0DEDB",x"10001",
									 x"0D6BA",x"10001",x"0DEBB",x"0D6BA",x"10001",x"0D69A",x"10002",x"0CE79",x"10002",x"0CE59",
									 x"10001",x"0C639",x"0C638",x"10001",x"0C618",x"0C639",x"0BDF7",x"09C90",x"07AE8",x"059E3",
									 x"05140",x"05980",x"061A0",x"06160",x"069C1",x"08282",x"0B463",x"0EE85",x"0FF05",x"0FEC5",
									 x"0FE44",x"0FE45",x"10000",x"0FE65",x"10000",x"0FE45",x"10000",x"0FE65",x"0FE45",x"10003",
									 x"0FE25",x"10002",x"0FE05",x"10000",x"0FDE5",x"0FDE4",x"0FDC4",x"0FDA4",x"10000",x"0FD84",
									 x"0FD63",x"0FD43",x"0FD04",x"0FCE4",x"0F4A3",x"0F462",x"0F463",x"0E4A8",x"0E590",x"0DE36",
									 x"0E6DA",x"0EF5D",x"0EF9E",x"0F7DF",x"0FFFF",x"10009",x"0FFFF",x"1000B",x"0F7BE",x"0EF7D",
									 x"0E71B",x"0DE98",x"0E614",x"0E50C",x"0EC45",x"0F463",x"0F483",x"0F4C3",x"0F503",x"0FD23",
									 x"0FD64",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"10000",x"0FDE5",x"0FE05",x"10000",x"0FE25",
									 x"10001",x"0FE45",x"10009",x"0FE65",x"10000",x"0FEA5",x"0FF06",x"0FF46",x"0D605",x"09382",
									 x"06180",x"05920",x"061A0",x"061C0",x"05980",x"04940",x"05A24",x"08BEC",x"0AD33",x"0CE38",
									 x"0C638",x"0C618",x"0C638",x"10000",x"0CE59",x"10000",x"0CE79",x"10002",x"0D69A",x"10001",
									 x"0D6BA",x"10002",x"0DEDB",x"10003",x"0DEFB",x"10004",x"0E71C",x"10000",x"0E73C",x"10000",
									 x"0E71C",x"10001",x"0E73C",x"10003",x"0E73D",x"0EF5D",x"0EF7D",x"10005",x"0F79D",x"0F79E",
									 x"10002",x"0F7BE",x"10005",x"0F7DE",x"10003",x"0F7BE",x"10004",x"0F79E",x"10001",x"0F79D",
									 x"0EF7D",x"10005",x"0EF5D",x"10001",x"0E75C",x"0E73C",x"10004",x"0E71C",x"10005",x"0DEFB",
									 x"10001",x"0DEDB",x"10003",x"0D6BA",x"10002",x"0D69A",x"10002",x"0CE79",x"10002",x"0CE59",
									 x"10000",x"0C638",x"0C618",x"0BE18",x"0C659",x"10000",x"0B5B6",x"083AC",x"051E4",x"04981",
									 x"051A1",x"061A0",x"06181",x"05940",x"07222",x"09363",x"0CD65",x"0F6C6",x"0FEE5",x"0FEA5",
									 x"0FE45",x"10001",x"0FE65",x"10000",x"0FE45",x"10000",x"0FE65",x"0FE45",x"10003",x"0FE25",
									 x"10002",x"0FE05",x"10000",x"0FDE5",x"0FDC4",x"10000",x"0FDA4",x"10000",x"0FD84",x"0FD63",
									 x"0FD23",x"0FD04",x"0F4C4",x"0F483",x"0F462",x"0F444",x"0E4EA",x"0DE14",x"0DE78",x"0E6DA",
									 x"0EF7D",x"0F7BE",x"0FFFF",x"1000A",x"0FFFF",x"1000B",x"0F7BE",x"0EF7D",x"0E71C",x"0DEBA",
									 x"0E677",x"0E54E",x"0E466",x"0F443",x"0F483",x"0F4C3",x"0F4E3",x"0F503",x"0FD43",x"0FD64",
									 x"0FD84",x"0FDA4",x"0FDC4",x"10000",x"0FDE5",x"0FDE4",x"0FE05",x"10001",x"0FE25",x"10001",
									 x"0FE45",x"10001",x"0FE65",x"0FE45",x"0FE65",x"10004",x"0F664",x"0FEE5",x"0FF46",x"0DE64",
									 x"09C01",x"061E0",x"05940",x"061A0",x"10000",x"05960",x"04920",x"051E3",x"07B6A",x"0A4B0",
									 x"0CE37",x"0C638",x"10002",x"0CE59",x"10000",x"0CE79",x"10001",x"0D69A",x"10002",x"0D6BA",
									 x"10002",x"0DEDB",x"10003",x"0DEFB",x"10002",x"0E71C",x"10000",x"0E73C",x"10004",x"0EF5D",
									 x"10006",x"0EF7D",x"10000",x"0F79E",x"10002",x"0EF7D",x"0F79E",x"10003",x"0F7BE",x"10004",
									 x"0F7DE",x"10008",x"0F7BE",x"10001",x"0F79E",x"10003",x"0EF7D",x"0F79E",x"10000",x"0EF7D",
									 x"10003",x"0EF5D",x"10001",x"0E75D",x"10000",x"0E73C",x"10004",x"0E71C",x"10002",x"0DEFB",
									 x"10001",x"0DEDB",x"10003",x"0D6BA",x"10002",x"0D69A",x"10001",x"0CE79",x"10002",x"0CE59",
									 x"0C638",x"10001",x"0C618",x"0C659",x"0C639",x"0AD34",x"07B4A",x"04981",x"04960",x"059C1",
									 x"061A0",x"06181",x"05100",x"07A61",x"0A3E2",x"0DDE5",x"0FF06",x"0FEA5",x"0FE85",x"0FE44",
									 x"0FE45",x"10000",x"0FE64",x"0FE45",x"10007",x"0FE24",x"0FE25",x"10000",x"0FE05",x"10000",
									 x"0FDE5",x"10000",x"0FDC4",x"0FDA4",x"0FD84",x"10000",x"0FD64",x"0FD63",x"0FD23",x"0FCE4",
									 x"0F4C3",x"0F483",x"0F463",x"0EC45",x"0E52D",x"0DE57",x"0D6BB",x"0E6FB",x"0EF7D",x"0F7BE",
									 x"0FFFF",x"1000A",x"0FFFF",x"1000B",x"0FFDF",x"0F79E",x"0E73D",x"0DEFC",x"0DE98",x"0DD91",
									 x"0E4A9",x"0EC44",x"0F463",x"0F4A3",x"0F4E3",x"0F503",x"0FD23",x"0FD64",x"0FD84",x"0FDA4",
									 x"10000",x"0FDC4",x"0FDE4",x"10000",x"0FE05",x"10001",x"0FE25",x"10001",x"0FE45",x"10001",
									 x"0FE65",x"0FE45",x"0FE65",x"10004",x"0F664",x"0FEC5",x"0FF26",x"0EEC4",x"0ACE1",x"07AA0",
									 x"069C1",x"06180",x"10000",x"05980",x"05140",x"04961",x"05A45",x"083AB",x"0BD95",x"0D679",
									 x"0CE79",x"0CE39",x"0C639",x"0C638",x"0CE59",x"10001",x"0CE79",x"0D69A",x"10002",x"0D6BA",
									 x"10002",x"0DEDB",x"10004",x"0DEFB",x"10001",x"0E71C",x"10000",x"0E73C",x"10003",x"0EF5D",
									 x"10001",x"0EF5C",x"0EF7D",x"10003",x"0F79E",x"10004",x"0F7BE",x"0F79E",x"10000",x"0F7BE",
									 x"0F7BF",x"10000",x"0F7BE",x"0F7DF",x"1000B",x"0F7BE",x"10002",x"0F7BF",x"10000",x"0F7BE",
									 x"10001",x"0F79E",x"10003",x"0EF7D",x"10005",x"0EF5D",x"10000",x"0EF3D",x"10000",x"0EF3C",
									 x"10000",x"0E73C",x"10001",x"0E71C",x"10001",x"0DEFB",x"10001",x"0DEDB",x"10003",x"0D6BA",
									 x"10002",x"0D69A",x"10001",x"0CE79",x"10002",x"0CE58",x"0C638",x"10000",x"0CE59",x"10000",
									 x"0CE39",x"0BDD6",x"0942E",x"05A04",x"04140",x"04960",x"059A1",x"061A0",x"06180",x"05940",
									 x"08B02",x"0B4A2",x"0E665",x"0FF26",x"0FEA5",x"0FE65",x"0FE45",x"10001",x"0FE64",x"0FE45",
									 x"10007",x"0FE24",x"10000",x"0FE25",x"0FE05",x"10000",x"0FDE5",x"0FDE4",x"0FDC4",x"0FDA4",
									 x"0FD84",x"10000",x"0FD64",x"0FD43",x"0F503",x"0FCE4",x"0F4A3",x"0F463",x"0EC64",x"0EC88",
									 x"0E570",x"0DE79",x"0DEFC",x"0E71C",x"0F79E",x"0FFDF",x"0FFFF",x"1000A",x"0FFFF",x"1000B",
									 x"0FFDF",x"0F7BE",x"0EF5D",x"0E71C",x"0DEBA",x"0E5F3",x"0ED0B",x"0EC65",x"0F463",x"0F4A3",
									 x"0F4C3",x"0F4E3",x"0F523",x"0FD44",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"10001",x"0FDE5",
									 x"0FE05",x"10000",x"0FE25",x"10001",x"0FE45",x"10001",x"0FE65",x"0FE45",x"0FE65",x"10000",
									 x"0FE85",x"0FE65",x"10002",x"0FEA5",x"0FF06",x"0F725",x"0CDC3",x"09BA2",x"07A42",x"06160",
									 x"06180",x"06181",x"05981",x"04960",x"04181",x"05A45",x"08C0E",x"0B596",x"0C618",x"0CE5A",
									 x"0D69A",x"0CE9A",x"0CE79",x"10002",x"0D69A",x"10001",x"0D6BA",x"10003",x"0DEDB",x"10002",
									 x"0DEFB",x"10003",x"0E71C",x"0E73C",x"10003",x"0EF5D",x"10003",x"0EF7D",x"10002",x"0F79D",
									 x"0F79E",x"10002",x"0F7BE",x"10000",x"0F7BF",x"10002",x"0F7DF",x"0FFDF",x"0FFFF",x"1000D",
									 x"0FFDF",x"10003",x"0F7DF",x"0F7BF",x"10001",x"0F7BE",x"10001",x"0F79E",x"10001",x"0EF9E",
									 x"0EF9D",x"0EF7D",x"10002",x"0EF5D",x"0EF3D",x"10000",x"0EF5D",x"0EF3D",x"0E73C",x"10001",
									 x"0E71C",x"10001",x"0DEFB",x"10002",x"0DEDB",x"10003",x"0D6BA",x"10001",x"0D69A",x"10002",
									 x"0CE79",x"10000",x"0CE59",x"0CE79",x"10000",x"0CE7A",x"0D67A",x"0CE18",x"0AD13",x"0942F",
									 x"06267",x"04140",x"04960",x"051A1",x"061C2",x"061A0",x"06180",x"061A0",x"0A3E4",x"0CDA4",
									 x"0EEA5",x"0FF06",x"0FE85",x"0FE45",x"10002",x"0FE64",x"0FE45",x"10007",x"0FE24",x"0FE04",
									 x"10001",x"0FDE4",x"10000",x"0FDC4",x"10000",x"0FDA4",x"0FD84",x"10000",x"0FD64",x"0F543",
									 x"0F503",x"0F4C3",x"0F482",x"0EC43",x"0E465",x"0E4EB",x"0E5D2",x"0DE99",x"0DF1C",x"0EF5D",
									 x"0F7BE",x"0FFDF",x"0FFFF",x"1000A",x"0FFFF",x"1000C",x"0F7BE",x"0F79D",x"0DF3C",x"0DEDB",
									 x"0DE16",x"0E56F",x"0E466",x"0F463",x"0F462",x"0FCC3",x"0FCE3",x"0F504",x"0FD44",x"0FD63",
									 x"0FD84",x"0FDA5",x"0FDC4",x"10000",x"0FDE5",x"0FE05",x"10001",x"0FE25",x"10000",x"0FE45",
									 x"10001",x"0FE65",x"10008",x"0FE85",x"0FEC6",x"0FF45",x"0E664",x"0AC62",x"082C3",x"05940",
									 x"06180",x"061C0",x"10000",x"05180",x"04960",x"04961",x"05A86",x"0944F",x"0AD53",x"0CE59",
									 x"0D6DB",x"10000",x"0D69A",x"0CE7A",x"0D69A",x"0CE99",x"0CE79",x"0CE99",x"0D699",x"0D69A",
									 x"0D6BA",x"0D69A",x"0DEDA",x"10000",x"0D6BA",x"0DEDB",x"10001",x"0DEFB",x"10002",x"0E71C",
									 x"10001",x"0E73C",x"10002",x"0EF5D",x"10002",x"0EF7D",x"10002",x"0F79E",x"10002",x"0F7BE",
									 x"10004",x"0FFDF",x"10004",x"0FFFF",x"1000C",x"0FFDF",x"10004",x"0F7BE",x"10004",x"0F79E",
									 x"10001",x"0EF7D",x"10002",x"0EF5D",x"10004",x"0E73C",x"10001",x"0E71C",x"10000",x"0DEFB",
									 x"10000",x"0E71C",x"0DEFC",x"0DEFB",x"10001",x"0DEDA",x"10000",x"0D6BA",x"10000",x"0D69A",
									 x"0D6BA",x"10000",x"0D699",x"0D6B9",x"0D699",x"0D69A",x"10000",x"0CE79",x"0CE7A",x"0D6BA",
									 x"0D6DA",x"0D679",x"0B594",x"07BAC",x"06287",x"04982",x"04140",x"05180",x"059A1",x"061A1",
									 x"06181",x"06981",x"07260",x"0B4C3",x"0E645",x"0F6E6",x"0FEC5",x"0FE64",x"0FE65",x"0FE45",
									 x"10001",x"0FE44",x"0FE64",x"0FE45",x"10004",x"0FE25",x"0FE24",x"0FE04",x"10001",x"0FE05",
									 x"0FDE5",x"10000",x"0FDC4",x"10000",x"0FDA4",x"0FD84",x"0FD64",x"0F563",x"0F523",x"0F4E2",
									 x"0FCC3",x"0F482",x"0F463",x"0EC46",x"0DD0E",x"0DE56",x"0DEB8",x"0E71B",x"0EF9D",x"0F7DF",
									 x"0FFDF",x"0FFFF",x"1000A",x"0FFFF",x"1000C",x"0FFDF",x"0F7BE",x"0E73C",x"0DEDB",x"0DE58",
									 x"0E591",x"0E4A8",x"0F464",x"0F463",x"0FCA2",x"0FCE3",x"0F504",x"0FD43",x"0FD63",x"0FD84",
									 x"0FDA4",x"0FDC5",x"0FDC4",x"0FDE5",x"10000",x"0FE05",x"10000",x"0FE25",x"10000",x"0FE45",
									 x"10001",x"0FE65",x"10008",x"0FE85",x"0FEA5",x"0FF46",x"0EEC5",x"0BD04",x"08B43",x"06180",
									 x"06160",x"061A0",x"061E0",x"059C0",x"04980",x"04160",x"051E3",x"06AE8",x"083AC",x"09CD1",
									 x"0B595",x"0BDD7",x"0CE59",x"0D6BB",x"0DEDB",x"10000",x"0D6DA",x"0D6BA",x"10001",x"0D6BB",
									 x"0DEDB",x"10000",x"0D6BB",x"0D6BA",x"0DEDB",x"10001",x"0DEFB",x"10002",x"0E71C",x"10000",
									 x"0E73C",x"10003",x"0EF5D",x"10002",x"0EF7D",x"10002",x"0F79E",x"10002",x"0F7BE",x"10004",
									 x"0FFDF",x"10004",x"0FFFF",x"1000C",x"0FFDF",x"10004",x"0F7BE",x"10004",x"0F79E",x"10001",
									 x"0EF7D",x"10002",x"0EF5D",x"10004",x"0E73C",x"10001",x"0E71C",x"10001",x"0DEFB",x"0DEFC",
									 x"10000",x"0DEFB",x"0DEDB",x"10000",x"0DEDA",x"10000",x"0D6DA",x"0D6BA",x"10000",x"0D69A",
									 x"0CE9A",x"0D6BA",x"10000",x"0D6DB",x"0DEDB",x"10000",x"0D6BA",x"0CE79",x"0BDF6",x"0B574",
									 x"0A4F2",x"08BED",x"05A66",x"051E3",x"04981",x"04960",x"051A0",x"061A1",x"10000",x"06160",
									 x"06981",x"082E0",x"0C564",x"0EEC6",x"0FEE6",x"0FEC4",x"0FE64",x"0FE44",x"0FE65",x"10001",
									 x"0FE64",x"0FE65",x"10001",x"0FE45",x"10002",x"0FE25",x"0FE24",x"0FE04",x"10001",x"0FE05",
									 x"0FDE4",x"10000",x"0FDC4",x"0FDA4",x"10000",x"0FD64",x"0FD44",x"0F543",x"0F523",x"0F4E2",
									 x"0FCC2",x"0F483",x"0F464",x"0E488",x"0DD70",x"0DE78",x"0DEBA",x"0E73C",x"0F79E",x"0FFDF",
									 x"0FFFF",x"1000B",x"0FFFF",x"1000D",x"0F7DF",x"0E77D",x"0DF1C",x"0E6DA",x"0E614",x"0DCEC",
									 x"0EC87",x"0EC44",x"0F482",x"0FCC2",x"0FCE3",x"0FD23",x"0FD63",x"0FD84",x"0FDA4",x"0FDA5",
									 x"0FDC4",x"10000",x"0FDE5",x"0FE05",x"10000",x"0FE25",x"10000",x"0FE45",x"10001",x"0FE65",
									 x"10009",x"0F685",x"0FF05",x"0F705",x"0D5E5",x"0AC65",x"07240",x"06180",x"061A1",x"069C1",
									 x"061E0",x"059A0",x"051A0",x"04940",x"04961",x"04182",x"05205",x"06AE9",x"0838C",x"09CB1",
									 x"0BDF6",x"0C617",x"0CE58",x"0D69A",x"0D6BA",x"0D6BB",x"0DEDC",x"0DEDB",x"10000",x"0DEBB",
									 x"10000",x"0DEDB",x"10002",x"0DEFB",x"0E71C",x"0DEFB",x"10000",x"0E71C",x"10000",x"0E73C",
									 x"10002",x"0EF5D",x"10003",x"0EF7D",x"10002",x"0F79E",x"10002",x"0F7BE",x"10004",x"0FFDF",
									 x"10004",x"0FFFF",x"1000C",x"0FFDF",x"10004",x"0F7BE",x"10004",x"0F79E",x"10001",x"0EF7D",
									 x"10002",x"0EF5D",x"10004",x"0E73C",x"10001",x"0E71C",x"10004",x"0DEFB",x"10001",x"0DEDB",
									 x"0DEFB",x"0D6DB",x"0DEDB",x"0DEDC",x"10000",x"0D6DC",x"10000",x"0D6BB",x"0D69A",x"0CE79",
									 x"0C637",x"0BDD6",x"0A512",x"083CD",x"062A8",x"05205",x"04182",x"04161",x"04160",x"05180",
									 x"059C0",x"061C0",x"061C1",x"069A1",x"06180",x"071E0",x"09BC2",x"0E666",x"0FF47",x"0FEE5",
									 x"0FE84",x"0FE44",x"10000",x"0FE65",x"10005",x"0FE45",x"10002",x"0FE25",x"0FE24",x"10000",
									 x"0FE04",x"10000",x"0FDE5",x"0FDE4",x"0FDC4",x"10000",x"0FDA4",x"0FD84",x"0FD64",x"0FD44",
									 x"0FD23",x"0F503",x"0F4C2",x"0FC82",x"0F463",x"0EC86",x"0E4CB",x"0E5D3",x"0E6DA",x"0E6FB",
									 x"0EF5D",x"0F7BE",x"0FFFF",x"1000C",x"0FFFF",x"1000E",x"0EF9E",x"0DF3D",x"0DEFB",x"0DE56",
									 x"0DD50",x"0E4CA",x"0EC45",x"0F483",x"0FCA2",x"0FCC3",x"0FD03",x"0F543",x"0FD64",x"0FD84",
									 x"0FDA4",x"0FDC4",x"10000",x"0FDE5",x"0FE05",x"10000",x"0FE25",x"10001",x"0FE45",x"10000",
									 x"0FE65",x"10003",x"0FE85",x"0FE65",x"0FE85",x"0FE65",x"10002",x"0FEC5",x"0FF05",x"0EEC6",
									 x"0CD65",x"08B01",x"069C1",x"06180",x"069E1",x"10000",x"061E0",x"059C0",x"05180",x"05160",
									 x"04960",x"04981",x"051C2",x"059E4",x"05205",x"062E9",x"0734B",x"083EE",x"0A4F2",x"0C617",
									 x"0D6BA",x"0E71C",x"10001",x"0E6FC",x"0DEFC",x"0DEDB",x"10000",x"0DEFB",x"10000",x"0E71C",
									 x"10001",x"0DEFB",x"0E71C",x"10000",x"0E73C",x"10002",x"0EF5D",x"10004",x"0EF7D",x"10001",
									 x"0F79E",x"10001",x"0F7BE",x"10005",x"0FFDF",x"10004",x"0FFFF",x"1000C",x"0FFDF",x"10004",
									 x"0F7BE",x"10004",x"0F79E",x"10003",x"0EF7D",x"10001",x"0EF5D",x"10003",x"0E73C",x"10000",
									 x"0E71C",x"10005",x"0DEFB",x"10001",x"0DEDB",x"0D6DB",x"0D6FB",x"0DEDB",x"0E6FC",x"10000",
									 x"0E71C",x"0DEDB",x"0C617",x"0A533",x"0842F",x"06B4B",x"062E8",x"05A66",x"051E4",x"049A3",
									 x"04982",x"04960",x"051A0",x"10000",x"059C0",x"06200",x"061E0",x"061A0",x"069A0",x"071E0",
									 x"082C1",x"0BCE4",x"0EEE6",x"0FF67",x"0FEE5",x"0FE64",x"0FE65",x"10000",x"0FE85",x"0FE65",
									 x"10004",x"0FE45",x"10002",x"0FE24",x"10000",x"0FE04",x"10000",x"0FDE4",x"10000",x"0FDC4",
									 x"10001",x"0FDA4",x"0FD84",x"0FD64",x"0FD23",x"0FD03",x"0F4E3",x"0F4A3",x"0F462",x"0EC44",
									 x"0E4C9",x"0DD4F",x"0DE36",x"0E6DB",x"0E71D",x"0EF7E",x"0FFDF",x"0FFFF",x"1000C",x"0FFFF",
									 x"1000D",x"0FFDF",x"0F79E",x"0E75D",x"0DF1B",x"0DE77",x"0DDB3",x"0E50D",x"0E466",x"0EC63",
									 x"0FC82",x"0FCA3",x"0FD04",x"0F543",x"0FD64",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FDE5",
									 x"0FE05",x"10000",x"0FE25",x"10001",x"0FE24",x"0FE45",x"0FE65",x"10003",x"0FE85",x"0FE65",
									 x"0FE85",x"10000",x"0FE65",x"10001",x"0FEA5",x"0FF05",x"0FF46",x"0DE46",x"09BE2",x"07200",
									 x"06180",x"069C0",x"06A01",x"10000",x"061C0",x"10000",x"059A0",x"051A0",x"04980",x"04140",
									 x"04940",x"04141",x"04182",x"049E4",x"05A66",x"07B6B",x"09C90",x"0AD53",x"0BDD5",x"0C5F6",
									 x"0CE58",x"0D699",x"0DEDB",x"0E71C",x"10000",x"0E73C",x"10002",x"0E71C",x"10002",x"0E73C",
									 x"10004",x"0EF5D",x"10002",x"0EF7D",x"10001",x"0F79E",x"10001",x"0F7BE",x"10005",x"0FFDF",
									 x"10004",x"0FFFF",x"1000C",x"0FFDF",x"10004",x"0F7BE",x"10004",x"0F79E",x"10003",x"0EF7D",
									 x"10001",x"0EF5D",x"10003",x"0E73C",x"10001",x"0E71C",x"10002",x"0E71B",x"10000",x"0E71C",
									 x"0E73C",x"0E71C",x"10001",x"0DEFB",x"0D69A",x"0CE38",x"0CE17",x"0BDD6",x"0B553",x"09CB0",
									 x"083AC",x"062A7",x"049E3",x"04181",x"04140",x"10000",x"04160",x"04960",x"04980",x"051C0",
									 x"059C0",x"061C0",x"061E0",x"069E0",x"069C0",x"10000",x"07220",x"09361",x"0CDC4",x"0F726",
									 x"0FF46",x"0FEC5",x"0FE45",x"10000",x"0FE65",x"0FE85",x"0FE65",x"10004",x"0FE45",x"10002",
									 x"0FE24",x"10000",x"0FE04",x"10000",x"0FDE4",x"10000",x"0FDC4",x"10000",x"0FDA4",x"10000",
									 x"0FD84",x"0FD43",x"0FD23",x"0FD03",x"0FCC3",x"0F483",x"0F462",x"0EC45",x"0E4EB",x"0D5B2",
									 x"0D657",x"0E6FB",x"0E73D",x"0EF7E",x"0FFDF",x"0FFFF",x"1000C",x"0FFFF",x"1000D",x"0FFDF",
									 x"0FFBE",x"0EF9E",x"0DF3C",x"0DE98",x"0DE16",x"0E54F",x"0E487",x"0EC63",x"0FC82",x"0FCA2",
									 x"0FD04",x"0F524",x"0FD43",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"10000",x"0FDE5",x"0FE05",
									 x"10000",x"0FE24",x"10001",x"0FE45",x"0FE65",x"10003",x"0FE85",x"0FE65",x"0FE85",x"10001",
									 x"0FE65",x"10000",x"0FE85",x"0FF04",x"0FF85",x"0EEC6",x"0B4A4",x"08261",x"069A0",x"069C0",
									 x"07201",x"10000",x"061C0",x"061E1",x"059E0",x"10000",x"051C0",x"051A0",x"04960",x"10000",
									 x"04140",x"10000",x"03961",x"041A2",x"049E3",x"05245",x"062A7",x"0734B",x"0946F",x"0AD54",
									 x"0CE59",x"0E71C",x"0E73C",x"1000A",x"0EF5D",x"10005",x"0EF7D",x"0EF9E",x"0F79E",x"10002",
									 x"0F7BE",x"10005",x"0FFDF",x"10004",x"0FFFF",x"1000C",x"0FFDF",x"10003",x"0F7DE",x"0F7BE",
									 x"10004",x"0F79E",x"10002",x"0F79D",x"0EF7D",x"10001",x"0EF5D",x"10003",x"0E73C",x"10008",
									 x"0EF5D",x"10000",x"0E73D",x"0E71C",x"0D679",x"0B555",x"08C2F",x"07B8C",x"062C8",x"05245",
									 x"049C4",x"04182",x"04161",x"04140",x"10001",x"04980",x"05180",x"051A0",x"059C1",x"059E0",
									 x"06201",x"06A01",x"10000",x"07201",x"061A0",x"069C0",x"08AC1",x"0AC62",x"0EEA6",x"0F745",
									 x"0F704",x"0FEA5",x"0FE46",x"0FE45",x"0FE65",x"0FE85",x"0FE64",x"0FE65",x"10003",x"0FE45",
									 x"10002",x"0FE24",x"10000",x"0FE04",x"10000",x"0FDE4",x"10001",x"0FDC4",x"0FDA4",x"0FD84",
									 x"0FD63",x"0FD43",x"0FD23",x"0FCE3",x"0FCA3",x"0F483",x"0F443",x"0EC66",x"0E52D",x"0D635",
									 x"0CE98",x"0E71B",x"0EF7D",x"0F7BE",x"0FFFF",x"1000D",x"0FFFF",x"1000E",x"0F7DF",x"0F7BE",
									 x"0E73C",x"0DEBA",x"0DE78",x"0DDD3",x"0DCEB",x"0EC66",x"0F443",x"0F483",x"0FCE4",x"0F503",
									 x"0FD23",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"10001",x"0FDE4",x"0FE05",x"0FE25",x"10000",
									 x"0FE45",x"0FE25",x"0FE45",x"10000",x"0FE65",x"10003",x"0FE85",x"10002",x"0FE65",x"0FE64",
									 x"0FEE4",x"0FF65",x"0FF26",x"0D5E4",x"09BA1",x"07A40",x"071C0",x"069C0",x"07200",x"07221",
									 x"07241",x"06A20",x"10000",x"06200",x"059E0",x"059C0",x"051A0",x"10000",x"04980",x"04160",
									 x"04140",x"03920",x"03120",x"03961",x"049C3",x"05245",x"062C8",x"07B6B",x"08C2E",x"09490",
									 x"0A4D1",x"0B574",x"0BDD6",x"0CE78",x"0DEDB",x"0E73C",x"0EF5D",x"0EF7D",x"10001",x"0EF7E",
									 x"10000",x"0EF7D",x"10005",x"0F77D",x"0F77E",x"0F79E",x"10001",x"0F7BE",x"10001",x"0FF9E",
									 x"0F79E",x"0FFBE",x"0FFDE",x"0FFDF",x"10003",x"0FFFF",x"1000C",x"0FFDF",x"10000",x"0FFDE",
									 x"10003",x"0F7BE",x"10001",x"0FFBE",x"0F7BE",x"10000",x"0F79E",x"10000",x"0F79D",x"0F79E",
									 x"0F79D",x"10000",x"0EF7D",x"10004",x"0EF5D",x"10000",x"0EF7D",x"10001",x"0EF9E",x"0EF5D",
									 x"0E73C",x"0DF1B",x"0CE78",x"0BDB6",x"0B554",x"0A4F2",x"09470",x"08C0E",x"07B8C",x"06AC8",
									 x"05225",x"049E3",x"03961",x"03120",x"10000",x"03940",x"04160",x"04980",x"10000",x"051A0",
									 x"059C0",x"059E1",x"061E1",x"06A01",x"07201",x"07221",x"10000",x"07A20",x"07A00",x"071C1",
									 x"07201",x"09BC2",x"0C582",x"0FF27",x"0FF26",x"0F6A4",x"0FE85",x"0FE65",x"10008",x"0FE45",
									 x"10002",x"0FE25",x"10001",x"0FE05",x"0FDE5",x"0FDC4",x"10000",x"0FDA4",x"10000",x"0FD84",
									 x"0FD43",x"0FD23",x"0FCE3",x"0FCC4",x"0F4A2",x"0EC82",x"0EC65",x"0E4AA",x"0DDB2",x"0D677",
									 x"0D6DA",x"0E73C",x"0F7BE",x"10000",x"0FFFF",x"1000D",x"0FFFF",x"1000E",x"0F7DF",x"0F7BF",
									 x"0EF5D",x"0E6DA",x"0DE99",x"0D615",x"0DD4E",x"0E487",x"0F443",x"0FC82",x"0FCE3",x"0F4E3",
									 x"0F523",x"0FD44",x"0FD84",x"0FDA4",x"0FDC4",x"10001",x"0FDE4",x"0FE05",x"0FE25",x"10002",
									 x"0FE45",x"10000",x"0FE65",x"10003",x"0FE85",x"10002",x"0FE65",x"10000",x"0FEC5",x"0FF25",
									 x"0FF66",x"0EEA6",x"0B4A3",x"08B21",x"07A01",x"071C0",x"07A01",x"07A21",x"07A41",x"07241",
									 x"07240",x"06A40",x"06A20",x"06221",x"06201",x"059E1",x"051C1",x"051A1",x"049A1",x"04981",
									 x"04160",x"10000",x"04161",x"03941",x"10001",x"04182",x"04A04",x"05A87",x"0734B",x"08C0E",
									 x"0A512",x"0C5D6",x"0D658",x"0DEBA",x"0DEDA",x"0DEFB",x"10000",x"0E71C",x"0E73C",x"0EF5D",
									 x"0EF7D",x"0F77D",x"0F79D",x"0F79E",x"10006",x"0F7BE",x"10001",x"0FFBF",x"0F7BF",x"0FFBE",
									 x"10000",x"0FFBF",x"10000",x"0FFDF",x"10000",x"0FFFF",x"1000D",x"0FFDF",x"10001",x"0FFDE",
									 x"0FFDF",x"10001",x"0FFDE",x"0F7BE",x"10007",x"0F79E",x"10003",x"0EF9E",x"0EF7D",x"0EF5D",
									 x"0EF5C",x"10000",x"0E73C",x"0E6FB",x"10000",x"0DEDA",x"0D699",x"0CE58",x"0C5F6",x"0A513",
									 x"08C0E",x"0734B",x"062A8",x"049E5",x"04183",x"03962",x"03941",x"03940",x"04160",x"04180",
									 x"10000",x"04980",x"049A0",x"051C0",x"10000",x"059E0",x"10000",x"06200",x"06A21",x"10000",
									 x"07221",x"07A21",x"10000",x"07A41",x"07A20",x"079E0",x"071E1",x"082A1",x"0B4C3",x"0D643",
									 x"0FF47",x"0FF06",x"0FEA5",x"0FE85",x"0FE65",x"10008",x"0FE45",x"10002",x"0FE25",x"10000",
									 x"0FE05",x"10000",x"0FDE5",x"0FDC4",x"10000",x"0FDA4",x"0FD84",x"0FD64",x"0FD43",x"0FD23",
									 x"0FCE3",x"0FCC4",x"0F482",x"0EC62",x"0EC66",x"0E50D",x"0DDF4",x"0D699",x"0D6FB",x"0E75C",
									 x"0F7BE",x"0FFDF",x"0FFFF",x"1000D",x"0FFFF",x"1000F",x"0FFDF",x"0F77D",x"0E71B",x"0DEB9",
									 x"0D657",x"0DDB1",x"0E4A9",x"0F443",x"0FC83",x"0FCC3",x"0F4E3",x"0F503",x"0FD44",x"0FD64",
									 x"0FD84",x"0FDA4",x"0FDC4",x"10000",x"0FDE4",x"0FE04",x"10000",x"0FE24",x"10000",x"0FE25",
									 x"0FE45",x"10000",x"0FE65",x"0FE85",x"10000",x"0FE65",x"10000",x"0FE85",x"10002",x"0FE65",
									 x"10000",x"0FEA5",x"0FEE4",x"0FF45",x"0F727",x"0C563",x"0A3E2",x"07A20",x"071A1",x"07A01",
									 x"08221",x"08261",x"10000",x"07A61",x"10000",x"07241",x"07221",x"06A21",x"06221",x"06200",
									 x"059E1",x"10000",x"051C0",x"051A0",x"10000",x"04980",x"04960",x"04140",x"04120",x"04140",
									 x"04181",x"04182",x"049E4",x"05A26",x"06288",x"06AC9",x"07B2B",x"0838C",x"08BEE",x"09490",
									 x"0A512",x"0AD54",x"0C617",x"0DEDA",x"0EF5C",x"0F79E",x"0FFDF",x"1000C",x"0F7DF",x"0FFDF",
									 x"10000",x"0FFFF",x"10017",x"0FFDF",x"10000",x"0F7DF",x"0FFFF",x"0F7DF",x"10002",x"0FFDF",
									 x"10006",x"0FFBE",x"0EF3C",x"0DEBA",x"0CE38",x"0B575",x"09CB2",x"09C70",x"08C2F",x"07B8C",
									 x"0732A",x"06B09",x"062A8",x"05226",x"051E4",x"049A3",x"04161",x"04140",x"10000",x"04160",
									 x"04980",x"10001",x"051A0",x"051C0",x"059E0",x"10000",x"06200",x"10000",x"06A20",x"06A40",
									 x"07241",x"10000",x"07A41",x"08241",x"08261",x"08241",x"07A00",x"071E0",x"07A20",x"09BA1",
									 x"0D5E4",x"0EEE5",x"0FF26",x"0FEE5",x"0FE85",x"10000",x"0FE65",x"10008",x"0FE45",x"10001",
									 x"0FE25",x"10000",x"0FE05",x"10000",x"0FDE5",x"0FDE4",x"0FDC4",x"0FDA4",x"0FD84",x"10000",
									 x"0FD64",x"0FD43",x"0FD03",x"0FCE3",x"0FCA3",x"0F483",x"0E463",x"0E487",x"0E570",x"0D636",
									 x"0D699",x"0DF1B",x"0EF7D",x"0FFBF",x"0FFDF",x"0FFFF",x"1000D",x"0FFFF",x"1000F",x"0FFDF",
									 x"0F79E",x"0EF5D",x"0DEDA",x"0D699",x"0DE15",x"0E50C",x"0F486",x"0F463",x"0F4A3",x"0F4C3",
									 x"0F4E3",x"0FD23",x"0FD64",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FDE4",x"0FE04",x"10000",
									 x"0FE24",x"0FE25",x"10000",x"0FE45",x"10000",x"0FE65",x"10000",x"0FE85",x"0FE65",x"10000",
									 x"0FE85",x"10000",x"0FE84",x"0FE85",x"10000",x"0FE66",x"0FE85",x"0FEA4",x"0FF05",x"0FF47",
									 x"0E685",x"0C544",x"09342",x"07A01",x"081E1",x"08221",x"08A61",x"08261",x"08281",x"10001",
									 x"07A61",x"10000",x"07261",x"07241",x"06A41",x"06221",x"06200",x"06201",x"061E1",x"059E0",
									 x"059C0",x"051A0",x"10001",x"04980",x"10000",x"04140",x"03920",x"03100",x"030E0",x"03900",
									 x"03941",x"04183",x"04A05",x"05A67",x"062C8",x"07B6B",x"0942E",x"0A4B1",x"0AD13",x"0B575",
									 x"0BDB6",x"0C5D6",x"0CE17",x"0CE37",x"0CE58",x"0D699",x"0DEFA",x"0E71B",x"0EF3C",x"0F77D",
									 x"0F79E",x"0FFDF",x"10000",x"0FFDE",x"0FFFF",x"1001B",x"0FFDF",x"0F7DE",x"0F7BE",x"0EF9D",
									 x"0EF5C",x"0E71B",x"0DEDA",x"0D69A",x"0D659",x"0CE38",x"0C617",x"0BDD6",x"0BD95",x"0B574",
									 x"0AD13",x"09CB0",x"08C0E",x"07B8C",x"06AE9",x"05A47",x"05205",x"041A3",x"03941",x"03100",
									 x"10000",x"03900",x"03920",x"04140",x"04960",x"04980",x"10000",x"051A0",x"059C0",x"059E0",
									 x"10000",x"06200",x"06220",x"06221",x"06A21",x"06A41",x"07241",x"07261",x"07A61",x"07A60",
									 x"07A81",x"08281",x"08261",x"08A61",x"08A81",x"08261",x"07A21",x"07A00",x"08AE1",x"0BCE3",
									 x"0EEC5",x"0FF66",x"0FF05",x"0FEA5",x"0FE85",x"0FE65",x"10009",x"0FE45",x"10001",x"0FE25",
									 x"0FE05",x"10000",x"0FDE5",x"10000",x"0FDC4",x"10000",x"0FDA4",x"0FD84",x"0FD64",x"0FD44",
									 x"0FD23",x"0F503",x"0F4C3",x"0FC83",x"0F484",x"0E486",x"0E4EB",x"0E5F3",x"0D678",x"0D6BA",
									 x"0E73C",x"0FFBE",x"0FFDF",x"0FFFF",x"1000E",x"0FFFF",x"10010",x"0FFDF",x"0EF7E",x"0DEDB",
									 x"0D6BB",x"0DE98",x"0DD90",x"0E4EA",x"0EC86",x"0F463",x"0F4A2",x"0F4E3",x"0FD03",x"0FD44",
									 x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",x"10000",x"0FE04",x"0FE24",x"10000",x"0FE25",
									 x"0FE45",x"10000",x"0FE65",x"10000",x"0FE85",x"0FE65",x"10000",x"0FE85",x"10000",x"0FE84",
									 x"0FE85",x"10000",x"0FE65",x"0FE66",x"0FE84",x"0FEC4",x"0FF26",x"0F746",x"0E686",x"0AC62",
									 x"08280",x"07A01",x"08220",x"08A61",x"08A81",x"10000",x"08AA1",x"10000",x"08A81",x"10000",
									 x"08281",x"08261",x"07A61",x"07261",x"10001",x"07241",x"06A41",x"10000",x"06200",x"10000",
									 x"059E0",x"10000",x"059E1",x"051C0",x"051A0",x"04980",x"10000",x"04960",x"10000",x"04160",
									 x"04140",x"03940",x"03941",x"03942",x"03921",x"03922",x"03942",x"041A4",x"05206",x"05A67",
									 x"06AE9",x"07B6B",x"083CD",x"0946F",x"0A4F2",x"0B554",x"0C5D6",x"0D638",x"0DEBA",x"0EF1B",
									 x"0F75C",x"0F79D",x"0F7BE",x"10001",x"0FFBE",x"10009",x"0FFDE",x"10004",x"0FFBE",x"10001",
									 x"0FFDE",x"0FFBE",x"10000",x"0F7BD",x"0F79D",x"10000",x"0F77D",x"0E71B",x"0DEB9",x"0D678",
									 x"0C616",x"0B574",x"0A4F2",x"09450",x"083ED",x"07B8C",x"06B0A",x"05AA8",x"049E5",x"041A3",
									 x"03942",x"03921",x"10000",x"03941",x"10000",x"04161",x"04141",x"04160",x"04180",x"04980",
									 x"10001",x"051A0",x"10000",x"059C0",x"059E0",x"06200",x"06201",x"06200",x"06220",x"10000",
									 x"06A41",x"07261",x"07260",x"10000",x"07A81",x"10000",x"082A1",x"10000",x"08AA1",x"10001",
									 x"08A81",x"08A61",x"08A62",x"08221",x"10000",x"082A1",x"0A422",x"0DE25",x"0F745",x"0FF66",
									 x"0FEE5",x"0FE85",x"0FE65",x"10000",x"0FE85",x"0FE65",x"10001",x"0FE85",x"0FE65",x"10000",
									 x"0FE85",x"0FE65",x"10000",x"0FE45",x"10001",x"0FE25",x"0FE05",x"10000",x"0FDE5",x"0FDC4",
									 x"10001",x"0FDA4",x"0FD84",x"0FD64",x"0FD44",x"0FD23",x"0F4E3",x"0F4A2",x"0F462",x"0EC45",
									 x"0E4CA",x"0DD6F",x"0E697",x"0DEDB",x"0D6FB",x"0EF5D",x"0FFDF",x"0FFFF",x"1000F",x"0FFFF",
									 x"10010",x"0FFDF",x"0F7BF",x"0DF1C",x"0D6FC",x"0D69A",x"0DDD3",x"0E52D",x"0E4A8",x"0EC63",
									 x"0FC82",x"0F4C3",x"0F503",x"0FD44",x"0FD64",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FDE4",
									 x"0FE04",x"0FE24",x"10001",x"0FE25",x"0FE45",x"0FE65",x"10000",x"0FE85",x"0FE65",x"10000",
									 x"0FE85",x"10000",x"0FE84",x"10000",x"0FEA4",x"0FE85",x"0FE66",x"0FE85",x"0FEA5",x"0FEE5",
									 x"0FF67",x"0EF06",x"0C543",x"09341",x"07A40",x"08220",x"08A41",x"09281",x"092A1",x"10003",
									 x"09281",x"08A81",x"10000",x"08281",x"07A81",x"10000",x"07260",x"07261",x"06A40",x"10001",
									 x"06220",x"06200",x"06220",x"05A00",x"059E0",x"051E0",x"059E0",x"051C0",x"051A0",x"05180",
									 x"04960",x"10000",x"04120",x"04100",x"03900",x"038E0",x"03100",x"03921",x"04161",x"04982",
									 x"051E4",x"05A25",x"05A67",x"06AA8",x"0732A",x"07B6B",x"083AD",x"08BEF",x"09450",x"09C71",
									 x"0A4B1",x"0A512",x"0AD33",x"0AD54",x"0B554",x"0B574",x"10000",x"0BD95",x"0BDB5",x"0BDB6",
									 x"0C5D6",x"0C5F6",x"0C5F7",x"0C617",x"0CE17",x"10003",x"0C617",x"0C5F7",x"0C5D6",x"0BDB6",
									 x"0BD95",x"0B575",x"0B574",x"10000",x"0B553",x"0AD33",x"0AD13",x"0A4F2",x"0A4D2",x"09C70",
									 x"0942F",x"08C0E",x"083CD",x"07B6B",x"0732A",x"06AE8",x"05A87",x"05245",x"04A04",x"041A2",
									 x"03941",x"03920",x"10000",x"03900",x"10000",x"03920",x"04140",x"04960",x"10000",x"051A0",
									 x"10000",x"051C0",x"10000",x"059C0",x"059E0",x"06200",x"06220",x"10000",x"06A40",x"06A41",
									 x"06A61",x"10000",x"07261",x"07281",x"10000",x"07A80",x"08280",x"082A1",x"10000",x"08AA1",
									 x"10002",x"092A1",x"09281",x"09282",x"08A42",x"08201",x"08241",x"09341",x"0BCE3",x"0EEE6",
									 x"0FF45",x"10000",x"0FEC4",x"0FE85",x"0FE65",x"0FE64",x"0FE84",x"0FE65",x"10007",x"0FE45",
									 x"10001",x"0FE25",x"0FE05",x"10000",x"0FDE5",x"0FDC4",x"10000",x"0FDA4",x"10000",x"0FD84",
									 x"0FD64",x"0FD44",x"0FD03",x"0FCE3",x"0FCA2",x"0F462",x"0E466",x"0E52E",x"0D5D3",x"0DE78",
									 x"0DEFC",x"0DF3D",x"0EF7D",x"0FFDF",x"0FFFF",x"1000F",x"0FFFF",x"10011",x"0F7BE",x"0EF5D",
									 x"0DF1C",x"0CEBA",x"0D616",x"0E5B2",x"0E4EB",x"0EC64",x"0FC62",x"0F4C3",x"0FCE3",x"0F523",
									 x"0F544",x"0F563",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",x"0FE05",x"10000",x"0FE25",x"10000",
									 x"0FE45",x"10001",x"0FE65",x"0FE85",x"10009",x"0FEA5",x"10000",x"0FF46",x"0F746",x"0DE85",
									 x"0AC83",x"08B01",x"08260",x"08240",x"08A61",x"092A2",x"092C1",x"10000",x"092C2",x"10000",
									 x"092C1",x"10002",x"08AA1",x"10000",x"082A1",x"08281",x"07A81",x"07A61",x"10000",x"07261",
									 x"10001",x"06A41",x"10000",x"06A21",x"06220",x"06200",x"05A00",x"059E0",x"10001",x"059C0",
									 x"051A0",x"10001",x"049A0",x"04980",x"10001",x"04160",x"04141",x"10000",x"03921",x"10000",
									 x"03101",x"03102",x"03902",x"03102",x"10000",x"03922",x"03942",x"04163",x"041A3",x"049C4",
									 x"10000",x"049E4",x"05205",x"05245",x"05A66",x"06287",x"062C8",x"06AC8",x"10000",x"06AE9",
									 x"10004",x"062C8",x"06288",x"05A67",x"05A46",x"05226",x"049E5",x"049C4",x"041C4",x"041A4",
									 x"03983",x"03943",x"03122",x"03102",x"10001",x"03122",x"03121",x"03101",x"03921",x"03941",
									 x"04141",x"04160",x"10000",x"04980",x"10000",x"049A0",x"10000",x"051A0",x"051C0",x"059C0",
									 x"059E0",x"10001",x"06200",x"06201",x"06221",x"06241",x"06A41",x"10000",x"07241",x"07261",
									 x"07A81",x"10002",x"08281",x"082A1",x"10000",x"08AA1",x"092C1",x"092E2",x"092C2",x"092C1",
									 x"09AC2",x"092C2",x"10000",x"092A2",x"092A1",x"08A61",x"08A41",x"08200",x"08AE0",x"0AC81",
									 x"0D624",x"0FF87",x"0FF25",x"0FEE5",x"0FEA5",x"10000",x"0FE85",x"10001",x"0FE65",x"10005",
									 x"0FE45",x"10003",x"0FE25",x"0FE04",x"10000",x"0FDE4",x"0FDC4",x"0FDA4",x"0FD84",x"0FD64",
									 x"10000",x"0FD44",x"0FD23",x"0FD03",x"0FCA3",x"0FC82",x"0EC63",x"0DCA9",x"0DD92",x"0DE35",
									 x"0D678",x"0DF1C",x"0EF5D",x"0F7BE",x"0FFDF",x"0FFFF",x"1000F",x"0FFFF",x"10012",x"0F79E",
									 x"0E75D",x"0D6DC",x"0D679",x"0E635",x"0E54F",x"0EC87",x"0F463",x"0F482",x"0FCC3",x"0FD03",
									 x"0FD43",x"0F563",x"0FD83",x"0FDA4",x"10000",x"0FDC4",x"0FDE5",x"0FE05",x"0FE25",x"10000",
									 x"0FE45",x"10001",x"0FE65",x"0FE85",x"10009",x"0FEA5",x"10000",x"0FF06",x"0F725",x"0F767",
									 x"0D606",x"0A403",x"08AC1",x"08220",x"08A62",x"09282",x"09AC1",x"09AE1",x"09AE2",x"09B02",
									 x"10000",x"09B01",x"09B02",x"10000",x"09AE2",x"092E1",x"10000",x"092C2",x"08AC2",x"10001",
									 x"082C2",x"10001",x"07AA2",x"10000",x"07A82",x"07281",x"07261",x"06A61",x"10000",x"06A41",
									 x"10000",x"06241",x"06221",x"10001",x"06201",x"05A01",x"059E0",x"10000",x"051C0",x"051A0",
									 x"051A1",x"049A1",x"10002",x"04161",x"10000",x"04140",x"10002",x"03940",x"10000",x"04160",
									 x"04161",x"10000",x"03961",x"04181",x"10000",x"04182",x"10003",x"041A2",x"10000",x"04182",
									 x"10001",x"04181",x"10001",x"04161",x"04160",x"03960",x"04160",x"10002",x"03961",x"03960",
									 x"04160",x"04181",x"10000",x"049A1",x"10001",x"051C1",x"051C0",x"051E0",x"059E0",x"05A00",
									 x"10001",x"05A20",x"06220",x"10000",x"06241",x"06A41",x"10001",x"07261",x"07262",x"07281",
									 x"10000",x"07A81",x"07AA2",x"082A2",x"10000",x"08AC2",x"10001",x"08AE2",x"092E2",x"10002",
									 x"09B02",x"10000",x"09AE2",x"0A2E2",x"0A302",x"10000",x"09AE1",x"09AC1",x"09AA1",x"08A60",
									 x"08240",x"08A61",x"0AC22",x"0DE25",x"0EF06",x"0FF87",x"0FF05",x"0FEC5",x"0FE85",x"10003",
									 x"0FE65",x"10005",x"0FE45",x"10002",x"0FE25",x"10000",x"0FE04",x"0FDE4",x"10000",x"0FDC4",
									 x"0FDA4",x"0FD83",x"0FD64",x"10000",x"0FD23",x"0FD02",x"0FCC3",x"0F483",x"0F463",x"0EC85",
									 x"0DD2D",x"0DE16",x"0D678",x"0DEBA",x"0E73C",x"0F79E",x"0FFDF",x"0FFFF",x"10010",x"0FFFF",
									 x"10012",x"0FFDF",x"0EF9E",x"0DEFC",x"0D69A",x"0D658",x"0DDB2",x"0E4C9",x"0F444",x"0F463",
									 x"0FCA3",x"0FCE3",x"0FD23",x"0F543",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE5",x"0FE05",
									 x"10000",x"0FE25",x"10001",x"0FE45",x"0FE65",x"10003",x"0FE85",x"10007",x"0FEE6",x"0F705",
									 x"0FFA7",x"0E6A6",x"0BD04",x"09B82",x"08240",x"08A62",x"09282",x"09AC2",x"0A2E1",x"10000",
									 x"0A301",x"10002",x"0A302",x"0A301",x"09AE1",x"09B01",x"09AE1",x"10001",x"092C1",x"092E1",
									 x"08AC1",x"10000",x"082C1",x"10000",x"082A1",x"07AA1",x"10000",x"07A81",x"07281",x"07261",
									 x"10001",x"06A61",x"06A41",x"10001",x"06241",x"10000",x"06220",x"10001",x"06200",x"05A00",
									 x"10001",x"05A01",x"10000",x"059E0",x"051E0",x"10000",x"051C0",x"051A0",x"049A0",x"10003",
									 x"04180",x"10001",x"04160",x"10007",x"04180",x"10001",x"04980",x"049A0",x"10001",x"049C0",
									 x"10001",x"051E0",x"10002",x"059E0",x"10001",x"05A00",x"10001",x"06220",x"10001",x"06240",
									 x"10001",x"06A60",x"10002",x"07281",x"10001",x"07A81",x"07AA1",x"10000",x"082A1",x"10000",
									 x"08AC1",x"10000",x"092C1",x"092C2",x"092E2",x"10001",x"09AE1",x"10000",x"09B01",x"0A302",
									 x"10001",x"0A301",x"10001",x"0A2E1",x"09AE1",x"09AC0",x"092A0",x"08A40",x"08241",x"08B02",
									 x"0C524",x"0EEC6",x"0F746",x"0FF46",x"0FEE5",x"0FEC5",x"0FE84",x"0FE85",x"10005",x"0FE65",
									 x"10002",x"0FE45",x"10001",x"0FE25",x"10000",x"0FE05",x"0FE04",x"0FDE4",x"0FDC4",x"0FDA4",
									 x"10000",x"0FD83",x"0FD44",x"10000",x"0FD23",x"0FD03",x"0FCC3",x"0F484",x"0EC64",x"0E4C8",
									 x"0DD91",x"0D658",x"0D69A",x"0DEFB",x"0EF5D",x"0F7BE",x"0FFDF",x"0FFFF",x"10010",x"0FFFF",
									 x"10012",x"0FFDF",x"0F79E",x"0EF3C",x"0DEBA",x"0CE59",x"0DDF5",x"0E50C",x"0EC66",x"0EC64",
									 x"0F484",x"0FCA3",x"0FD03",x"0FD23",x"0FD64",x"10000",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE5",
									 x"0FE05",x"10000",x"0FE25",x"10000",x"0FE45",x"0FE65",x"10001",x"0FE85",x"10000",x"0FE65",
									 x"10000",x"0FE85",x"10005",x"0FEC6",x"0FF05",x"0FF65",x"0FF45",x"0E645",x"0BCC4",x"092E0",
									 x"08240",x"08A61",x"09AC2",x"0A2E1",x"0A2E0",x"0AB01",x"0AB21",x"0AB22",x"0AB21",x"10003",
									 x"0AB22",x"0A321",x"0A301",x"10000",x"09B01",x"10000",x"09301",x"10000",x"092E1",x"10000",
									 x"08AE1",x"08AC1",x"10000",x"082C1",x"082A1",x"10001",x"07AA1",x"07A81",x"10000",x"07281",
									 x"10000",x"07261",x"07241",x"10000",x"06A40",x"10002",x"06A41",x"10001",x"06221",x"06220",
									 x"06200",x"10001",x"05A00",x"10004",x"059E0",x"10000",x"059E1",x"10000",x"059E0",x"059C0",
									 x"10000",x"059E0",x"10000",x"059C0",x"059E0",x"10002",x"05A00",x"10004",x"05A20",x"06220",
									 x"10003",x"06A20",x"10000",x"06A40",x"06A60",x"10000",x"06A40",x"10000",x"07240",x"07261",
									 x"07281",x"10001",x"07A81",x"10000",x"07AA1",x"07AA0",x"082C1",x"10000",x"082E1",x"08AE1",
									 x"10000",x"092C1",x"092E1",x"09AE1",x"10000",x"09B01",x"0A301",x"0A302",x"10000",x"0A322",
									 x"10000",x"0A321",x"10000",x"0AB22",x"10000",x"0AB21",x"10000",x"0AB22",x"0A302",x"0A2E2",
									 x"10000",x"09AC1",x"09281",x"08A61",x"08AC2",x"0A423",x"0DE46",x"0F766",x"0FF66",x"0FF05",
									 x"0FEC5",x"0FEA5",x"10000",x"0FE85",x"10005",x"0FE65",x"10002",x"0FE45",x"10001",x"0FE25",
									 x"10000",x"0FE05",x"0FDE4",x"0FDC4",x"10000",x"0FDA4",x"0FD84",x"10000",x"0FD44",x"0FD24",
									 x"0FD03",x"0FCE3",x"0F484",x"0F464",x"0EC66",x"0DCEB",x"0DDF3",x"0D658",x"0D69A",x"0E71C",
									 x"0F79D",x"0FFDF",x"0FFFF",x"10011",x"0FFFF",x"10013",x"0FFDF",x"0F77D",x"0DEDB",x"0D69A",
									 x"0DE57",x"0E590",x"0E4CA",x"0ECA7",x"0EC65",x"0FC83",x"0FCC2",x"0FD23",x"0F544",x"0FD44",
									 x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE5",x"0FE05",x"0FE25",x"10000",x"0FE45",x"0FE65",
									 x"10002",x"0FE85",x"0FE65",x"0FE85",x"10006",x"0FEA5",x"0FEC5",x"0FF05",x"0FF65",x"0FF47",
									 x"0DE26",x"0B443",x"08AC0",x"08261",x"092A1",x"0A2E1",x"10000",x"0AB01",x"0AB21",x"0AB42",
									 x"10000",x"0AB62",x"10000",x"0B342",x"10001",x"0AB42",x"10001",x"0AB41",x"0A341",x"10000",
									 x"0A322",x"10001",x"09B22",x"09B21",x"10000",x"09301",x"10000",x"092E1",x"08AE1",x"10000",
									 x"08AC1",x"10000",x"082C1",x"10001",x"082C2",x"082A2",x"10001",x"07AA1",x"10000",x"07A81",
									 x"10000",x"07281",x"10001",x"07261",x"07262",x"07261",x"10000",x"06A61",x"10001",x"07261",
									 x"06A61",x"10004",x"06A41",x"10004",x"06A62",x"10000",x"06A61",x"10005",x"07282",x"10000",
									 x"07281",x"07A81",x"10005",x"07AA1",x"10000",x"082C2",x"10002",x"08AC2",x"08AE2",x"10001",
									 x"08AE1",x"092E1",x"09301",x"10000",x"09B21",x"09B22",x"10000",x"0A301",x"0A322",x"10000",
									 x"0AB22",x"0AB42",x"10004",x"0B341",x"10000",x"0AB42",x"10001",x"0AB22",x"10001",x"0A2E2",
									 x"10000",x"09282",x"08A60",x"09302",x"09BC2",x"0D5E6",x"0F747",x"0FF66",x"0FF46",x"0FEC5",
									 x"0FEA5",x"0FE84",x"0FE85",x"10006",x"0FE65",x"10002",x"0FE45",x"10000",x"0FE25",x"10001",
									 x"0FE05",x"0FDE4",x"0FDC4",x"0FDA4",x"0FD84",x"10000",x"0FD63",x"0FD24",x"0FD03",x"0FCE2",
									 x"0F4A2",x"0F463",x"0EC86",x"0E4CA",x"0E570",x"0DE56",x"0D699",x"0DEBA",x"0EF5D",x"0F7BE",
									 x"0FFFF",x"10012",x"0FFFF",x"10014",x"0F7BE",x"0E73C",x"0D6DB",x"0D6B9",x"0D615",x"0DD4F",
									 x"0E4CA",x"0EC66",x"0F463",x"0FCA2",x"0FD03",x"0F524",x"0FD44",x"0FD64",x"0FD84",x"0FDA4",
									 x"0FDC4",x"0FDE5",x"0FE05",x"10000",x"0FE24",x"10000",x"0FE45",x"0FE65",x"10001",x"0FE85",
									 x"10005",x"0FEA5",x"10003",x"0F6E5",x"0FF45",x"0FF86",x"0EEC6",x"0CD44",x"09340",x"08AC1",
									 x"08A81",x"09AC1",x"0A302",x"10000",x"0AB21",x"0AB22",x"0AB42",x"0AB62",x"0B362",x"10006",
									 x"0AB62",x"0AB42",x"10002",x"0A342",x"0A341",x"0A321",x"0A341",x"0A342",x"09B21",x"10000",
									 x"09B01",x"10000",x"09B02",x"09302",x"092E1",x"10000",x"08AE1",x"10001",x"08AE2",x"08AC1",
									 x"082C1",x"10003",x"082A1",x"07AA1",x"082C2",x"07AC1",x"07AA1",x"10003",x"07A81",x"07281",
									 x"10001",x"07A81",x"10000",x"07A61",x"07A81",x"10002",x"07281",x"07A81",x"10001",x"07AA1",
									 x"10007",x"07AC1",x"082C1",x"10002",x"082C2",x"082E2",x"08AE2",x"08AE1",x"10001",x"09301",
									 x"10002",x"09B01",x"10001",x"09B02",x"09B22",x"0A322",x"10002",x"0AB42",x"10003",x"0AB62",
									 x"10001",x"0B362",x"0B361",x"10001",x"0B362",x"10000",x"0AB62",x"0AB42",x"0A322",x"10000",
									 x"0A2E1",x"09AC2",x"08A81",x"08AA0",x"0A3C1",x"0B4C2",x"0EF06",x"0FFA7",x"0FF45",x"0FEE5",
									 x"0FEA5",x"10000",x"0FE85",x"0FEA5",x"10001",x"0FE85",x"10003",x"0FE65",x"10002",x"0FE45",
									 x"10000",x"0FE25",x"10000",x"0FE05",x"0FDE5",x"0FDC4",x"10000",x"0FDA4",x"0FD84",x"0FD64",
									 x"0FD44",x"0FD24",x"0FD03",x"0FCC2",x"0F4A2",x"0EC64",x"0E4C9",x"0DD2E",x"0DDD5",x"0D699",
									 x"0D6DA",x"0E6DB",x"0FFBE",x"0FFFF",x"10013",x"0FFFF",x"10014",x"0F7DF",x"0E77D",x"0DEFC",
									 x"0D6BA",x"0D637",x"0D5B2",x"0DD2C",x"0EC86",x"0F463",x"0F4A2",x"0FCE3",x"0FD23",x"0FD24",
									 x"0FD44",x"0FD84",x"0FDA4",x"0FDC4",x"10000",x"0FDE4",x"0FE05",x"0FE25",x"10000",x"0FE45",
									 x"10000",x"0FE65",x"10000",x"0FE85",x"10004",x"0FEA5",x"10000",x"0FE85",x"0FEA5",x"10001",
									 x"0FEC5",x"0FF05",x"0FF66",x"0F746",x"0DE65",x"0A440",x"09B62",x"08AA1",x"092A1",x"09AE1",
									 x"0A302",x"0AB22",x"0AB42",x"0AB62",x"0B362",x"0B382",x"10001",x"0B362",x"10000",x"0BB62",
									 x"0BB82",x"0B362",x"10002",x"0AB62",x"10000",x"0AB61",x"10000",x"0AB41",x"0AB42",x"10000",
									 x"0A322",x"0A321",x"09B21",x"10000",x"09B22",x"10001",x"09B01",x"10001",x"09301",x"10001",
									 x"092E1",x"08B02",x"10000",x"08AE2",x"10000",x"08AE1",x"08AC1",x"08AC2",x"10000",x"082C2",
									 x"10003",x"082C1",x"082C2",x"082A2",x"10000",x"082A1",x"10007",x"082C2",x"082C1",x"10004",
									 x"082C2",x"10001",x"08AC2",x"08AE2",x"08AE1",x"08AE2",x"10000",x"092E2",x"09302",x"10004",
									 x"09B21",x"10003",x"0A341",x"10000",x"0A342",x"10000",x"0AB42",x"10001",x"0AB62",x"10000",
									 x"0AB42",x"0B362",x"10003",x"0B382",x"10000",x"0BB82",x"0B382",x"10001",x"0B362",x"0B342",
									 x"0AB42",x"0AB22",x"0A302",x"09AE1",x"092A1",x"08A81",x"09341",x"0BCE3",x"0D624",x"0F786",
									 x"0FF66",x"0FF05",x"0FEA5",x"10003",x"0FE85",x"10003",x"0FE65",x"10004",x"0FE44",x"0FE45",
									 x"0FE25",x"0FE05",x"10000",x"0FDE5",x"0FDC4",x"0FDA4",x"10000",x"0FD84",x"0FD64",x"0FD23",
									 x"0FD03",x"0FCE3",x"0F4A2",x"0EC82",x"0E484",x"0E50C",x"0DDB2",x"0D616",x"0D699",x"0DEFB",
									 x"0E73C",x"0FFDF",x"0FFFF",x"10013",x"0FFFF",x"10015",x"0F7BF",x"0E75D",x"0DEDB",x"0D658",
									 x"0D616",x"0DD90",x"0E4C9",x"0EC64",x"0F483",x"0F4C3",x"0FD03",x"0FD23",x"0FD44",x"0FD64",
									 x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",x"0FE04",x"0FE05",x"0FE25",x"0FE45",x"10001",x"0FE65",
									 x"10000",x"0FE85",x"10004",x"0FEA5",x"0FE85",x"0FEA5",x"10001",x"0FEC5",x"0FEE5",x"0F705",
									 x"0FF66",x"0F746",x"0D604",x"0BCE5",x"09B42",x"092A1",x"092A0",x"0A2E2",x"0AB22",x"0AB42",
									 x"0AB41",x"0AB61",x"0B382",x"10000",x"0BB82",x"10006",x"0B3A2",x"10002",x"0B382",x"10001",
									 x"0B362",x"0AB62",x"10005",x"0A342",x"10005",x"09B42",x"10000",x"09B22",x"10003",x"09302",
									 x"10003",x"09322",x"09302",x"10001",x"09301",x"10006",x"09302",x"10000",x"09322",x"09302",
									 x"10001",x"09322",x"09302",x"09322",x"10002",x"09B22",x"10003",x"0A322",x"09B42",x"10000",
									 x"0A342",x"10003",x"0AB42",x"10000",x"0AB62",x"10002",x"0AB82",x"0B382",x"0B383",x"0B382",
									 x"10003",x"0BB82",x"10003",x"0BBA2",x"10001",x"0BB82",x"0B382",x"10000",x"0B362",x"10000",
									 x"0AB42",x"0AB22",x"0A2E2",x"092A1",x"08AA1",x"09301",x"0B4A4",x"0E687",x"0FF88",x"0FFA6",
									 x"0FF05",x"0FEC5",x"0FEA5",x"10003",x"0FE85",x"10002",x"0FE65",x"10004",x"0FE45",x"0FE44",
									 x"0FE24",x"0FE25",x"0FE05",x"0FDE5",x"0FDC5",x"0FDC4",x"0FDA4",x"0FD84",x"0FD64",x"10000",
									 x"0FD24",x"0FD04",x"0FCC3",x"0FC83",x"0EC64",x"0E4A8",x"0E56F",x"0DE15",x"0D678",x"0D6BA",
									 x"0EF5C",x"0EF9D",x"0FFFF",x"10014",x"0FFFF",x"10014",x"0FFFE",x"0FFFF",x"0F7BE",x"0E71C",
									 x"0DE79",x"0D658",x"0D5F4",x"0DD2D",x"0EC66",x"0F463",x"0F483",x"0FCC3",x"0F4E3",x"0FD23",
									 x"0FD44",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FDE4",x"0FE04",x"0FE05",x"0FE25",x"10000",
									 x"0FE45",x"0FE65",x"10002",x"0FE85",x"10002",x"0FEA5",x"0FE85",x"0FEA5",x"0FEC5",x"0FEA5",
									 x"0FEC5",x"10000",x"0F6E5",x"0FF46",x"0FF86",x"0FF67",x"0E686",x"0B483",x"092E0",x"08A81",
									 x"092A1",x"0A302",x"0AB42",x"0AB41",x"0AB61",x"0B382",x"0B3A2",x"0BBA2",x"10002",x"0C3A2",
									 x"0C3C2",x"0C3A2",x"0BBA2",x"0BBC2",x"0BBA2",x"0BBC2",x"0BBA2",x"0BBA1",x"0BBA2",x"10000",
									 x"0B3A2",x"0B382",x"10002",x"0B3A2",x"0B382",x"10001",x"0AB82",x"10002",x"0AB62",x"10000",
									 x"0AB61",x"10001",x"0AB41",x"10001",x"0A362",x"0A341",x"10003",x"0A361",x"09B41",x"1000F",
									 x"0A341",x"10006",x"0A361",x"0AB61",x"10003",x"0AB81",x"10001",x"0B381",x"0B382",x"0B383",
									 x"0B382",x"10003",x"0B3A2",x"0BBA2",x"1000D",x"0BB82",x"0B382",x"0B383",x"0B362",x"0AB42",
									 x"0AB21",x"0A301",x"092A1",x"08A81",x"09321",x"0A421",x"0DE46",x"0F747",x"0FFA7",x"0F725",
									 x"0FF05",x"0FEC5",x"0FEA5",x"10004",x"0FE85",x"10001",x"0FE65",x"10002",x"0FE45",x"10001",
									 x"0FE24",x"0FE25",x"0FE05",x"10000",x"0FDE5",x"0FDC4",x"0FDA4",x"0FD84",x"0FD64",x"0FD43",
									 x"0FD23",x"0F504",x"0F4C3",x"0FC83",x"0F463",x"0EC67",x"0E50D",x"0DDF3",x"0D657",x"0D6BA",
									 x"0DEFB",x"0F79D",x"0FFBE",x"0FFFF",x"10014",x"0FFFF",x"10016",x"0FFDF",x"0EF5D",x"0DEDB",
									 x"0D679",x"0CE57",x"0DDB1",x"0E4C9",x"0F464",x"0F463",x"0F4A3",x"0F4C3",x"0FD03",x"0FD24",
									 x"0FD64",x"0FDA4",x"10000",x"0FDC4",x"10000",x"0FDE4",x"0FE05",x"0FE25",x"10000",x"0FE45",
									 x"10000",x"0FE65",x"10002",x"0FE85",x"10001",x"0FEA5",x"10003",x"0FEC5",x"10000",x"0FEE5",
									 x"0FF26",x"0FF85",x"0FFA6",x"0F746",x"0DE05",x"0A401",x"09301",x"092C1",x"092E1",x"0A302",
									 x"0A321",x"0AB41",x"0B381",x"0B382",x"0BBA2",x"10002",x"0C3C2",x"10005",x"0BBC2",x"10004",
									 x"0BBA2",x"10006",x"0B3A2",x"10000",x"0B382",x"10005",x"0B362",x"0AB82",x"0AB62",x"10004",
									 x"0AB82",x"0AB62",x"10000",x"0A362",x"10004",x"0AB62",x"10001",x"0A362",x"10003",x"0AB62",
									 x"10008",x"0B362",x"0B382",x"10004",x"0BBA2",x"10008",x"0BBC2",x"10000",x"0C3C2",x"10001",
									 x"0BBC2",x"10000",x"0C3C2",x"10000",x"0BBC2",x"0BBA2",x"10003",x"0BB82",x"0B382",x"0B362",
									 x"0AB42",x"0AB22",x"0A301",x"09AE1",x"08AA0",x"09302",x"0AC22",x"0C563",x"0F726",x"0FF86",
									 x"0FF66",x"0FF05",x"0FEE5",x"0FEA5",x"10005",x"0FE85",x"10000",x"0FE65",x"10003",x"0FE45",
									 x"10001",x"0FE25",x"0FE04",x"0FE05",x"0FDE5",x"0FDC5",x"0FDA4",x"10000",x"0FD84",x"0FD44",
									 x"0FD23",x"10000",x"0F4E3",x"0F4C3",x"0F462",x"0F464",x"0E4C9",x"0DD91",x"0D636",x"0CE79",
									 x"0D6DC",x"0E75D",x"0FFBE",x"0FFDF",x"0FFFF",x"10014",x"0FFFF",x"10017",x"0F79E",x"0E6FC",
									 x"0D69A",x"0CE98",x"0D615",x"0DD2E",x"0EC87",x"0EC63",x"0F483",x"0F4A3",x"0FCE3",x"0FD23",
									 x"0FD44",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FDE4",x"0FDE5",x"0FE05",x"0FE25",x"10000",
									 x"0FE45",x"10002",x"0FE65",x"0FE85",x"10001",x"0FEA5",x"10003",x"0FEC5",x"10001",x"0FEE5",
									 x"0FF45",x"0FFA6",x"0FF86",x"0F727",x"0BD02",x"09BC1",x"09300",x"08AC0",x"09AE1",x"0A322",
									 x"0AB42",x"0AB62",x"0B382",x"10000",x"0BBA2",x"10001",x"0BBC2",x"0C3C2",x"1000A",x"0BBC2",
									 x"10007",x"0BBA2",x"10002",x"0B3A2",x"10005",x"0B382",x"1001E",x"0BB82",x"10000",x"0BB83",
									 x"10000",x"0BBA3",x"10001",x"0BBA2",x"10000",x"0BBA3",x"0C3C3",x"0C3C2",x"10003",x"0BBC2",
									 x"0C3C2",x"10006",x"0C3E2",x"0C3C2",x"0BBC2",x"10002",x"0BBA2",x"0B382",x"10000",x"0AB62",
									 x"0AB42",x"0A302",x"09AE1",x"092C0",x"08AE0",x"09BE1",x"0C564",x"0DE85",x"0FF66",x"0FF45",
									 x"0FF25",x"0FEE5",x"0FEE6",x"0FEA6",x"10000",x"0FEA5",x"0FEC5",x"0FEA5",x"10001",x"0FE85",
									 x"10001",x"0FE65",x"10002",x"0FE45",x"10000",x"0FE25",x"10000",x"0FE05",x"0FDE5",x"10000",
									 x"0FDC5",x"0FDA4",x"0FD84",x"0FD64",x"0FD44",x"0FD03",x"10000",x"0FCC2",x"0F4A3",x"0EC83",
									 x"0ECA7",x"0DD0D",x"0D5F5",x"0D679",x"0CE9A",x"0DF1D",x"0F79E",x"0FFBF",x"0FFDF",x"0FFFF",
									 x"10014",x"0FFFF",x"10017",x"0FFDF",x"0E75D",x"0DEDB",x"0D699",x"0CE17",x"0D592",x"0E4EB",
									 x"0EC65",x"0F464",x"0F482",x"0F4C3",x"0FD03",x"0FD23",x"0FD43",x"0FD84",x"0FDA4",x"10000",
									 x"0FDC4",x"0FDE5",x"0FE05",x"0FE25",x"10000",x"0FE45",x"10002",x"0FE65",x"0FE85",x"10001",
									 x"0FEA5",x"10003",x"0FEC5",x"10000",x"0FEA5",x"0FEC5",x"0FEE5",x"0FF46",x"0FF86",x"0FF87",
									 x"0E685",x"0CDA4",x"0AC02",x"09301",x"092C0",x"09AC1",x"0AB22",x"0AB62",x"10000",x"0B382",
									 x"10000",x"0BBA2",x"10000",x"0BBC2",x"10000",x"0C3E2",x"1000F",x"0C3E3",x"10000",x"0BBE3",
									 x"10000",x"0BBC3",x"10000",x"0BBC2",x"1000C",x"0BBA2",x"0BBC2",x"10003",x"0BBA2",x"10008",
									 x"0BBC2",x"10003",x"0BBA2",x"10000",x"0BBC2",x"10008",x"0C3C2",x"10003",x"0C3E2",x"10008",
									 x"0C3C2",x"10000",x"0C3E2",x"10001",x"0BBC2",x"10002",x"0BBA2",x"0B382",x"0B381",x"0AB62",
									 x"0AB22",x"09AE1",x"092C1",x"092E1",x"09BA1",x"0C563",x"0E6C7",x"0F767",x"0FF66",x"0FF06",
									 x"0FEE5",x"0FEC5",x"0FEC6",x"0FEA6",x"10000",x"0FEA5",x"0FEC5",x"0FEA5",x"10001",x"0FE85",
									 x"10001",x"0FE65",x"10002",x"0FE45",x"10000",x"0FE25",x"0FE05",x"10000",x"0FDE5",x"0FDC5",
									 x"0FDA4",x"10000",x"0FD84",x"0FD44",x"0FD23",x"0FCE3",x"10000",x"0F4A2",x"0EC84",x"0E4A6",
									 x"0E50B",x"0DD91",x"0D617",x"0DE9A",x"0DEDB",x"0E75E",x"0F7BF",x"0FFFF",x"10016",x"0FFFF",
									 x"10018",x"0F79E",x"0E73C",x"0DEDB",x"0D659",x"0D5F6",x"0DD50",x"0E4CA",x"0EC85",x"0F483",
									 x"0F4A2",x"0FCE2",x"0FD03",x"0FD24",x"0F564",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",x"0FE04",
									 x"0FE05",x"0FE04",x"0FE25",x"0FE45",x"10001",x"0FE65",x"10000",x"0FE85",x"10000",x"0FEA5",
									 x"10000",x"0FE85",x"0FEA5",x"10003",x"0FEC5",x"0FEE5",x"0FF05",x"0FF46",x"0FF67",x"0FF47",
									 x"0EEE6",x"0CD64",x"0A3E1",x"09300",x"092E1",x"09B02",x"0AB62",x"10001",x"0B382",x"0B3A2",
									 x"0BBC3",x"10000",x"0BBE3",x"0BBE2",x"0C3E2",x"10003",x"0C3E3",x"10001",x"0C3E2",x"10004",
									 x"0C3E3",x"10003",x"0C3E2",x"10004",x"0C3C2",x"10001",x"0C3E2",x"10001",x"0BBE2",x"10002",
									 x"0C3C2",x"10001",x"0C3E2",x"10000",x"0C3C2",x"0C3C3",x"10003",x"0C3C2",x"10004",x"0C3E2",
									 x"0BBC2",x"10004",x"0BBE2",x"0C3E2",x"1000F",x"0C3E3",x"0C403",x"10000",x"0C3E2",x"10006",
									 x"0BBE2",x"0BBC2",x"10002",x"0B3A2",x"0B381",x"0AB41",x"0A322",x"0A302",x"092C1",x"09301",
									 x"0A3A1",x"0BCE3",x"0E6A5",x"0FF68",x"0FF87",x"0FF26",x"0FEE6",x"0FEC5",x"0FEA5",x"10000",
									 x"0FEC5",x"10002",x"0FEA5",x"10001",x"0FE85",x"10002",x"0FE65",x"10000",x"0FE45",x"10000",
									 x"0FE25",x"0FE24",x"0FE04",x"0FDE4",x"10000",x"0FDC4",x"0FDA4",x"0FD64",x"10000",x"0F543",
									 x"0FD03",x"0FCE2",x"0F4A3",x"0F462",x"0EC85",x"0E4C9",x"0DD4F",x"0DDF4",x"0CE59",x"0D6BB",
									 x"0E73C",x"0EF9E",x"0FFDF",x"0FFFF",x"10016",x"0FFFF",x"10018",x"0F7BE",x"0EF9E",x"0E73C",
									 x"0D699",x"0D657",x"0D5D3",x"0DD2E",x"0E4A8",x"0EC64",x"0F482",x"0FCA2",x"0FCE3",x"0FD24",
									 x"0FD44",x"0FD84",x"10000",x"0FDA4",x"0FDC4",x"0FDE4",x"0FE04",x"10000",x"0FE25",x"0FE45",
									 x"10000",x"0FE65",x"10002",x"0FE85",x"10000",x"0FEA5",x"0FE85",x"0FEA5",x"10002",x"0FEC5",
									 x"10000",x"0FEE5",x"10000",x"0FF05",x"0FF46",x"0FF87",x"0FF88",x"0E686",x"0BD03",x"09360",
									 x"09301",x"092E1",x"0A322",x"0AB62",x"10000",x"0B382",x"10000",x"0B3A2",x"0B3C3",x"0BBC3",
									 x"0BBE2",x"10000",x"0C3E2",x"10002",x"0C3E3",x"10000",x"0C403",x"0C402",x"10000",x"0C3E2",
									 x"10000",x"0C402",x"0C3E2",x"0C3E3",x"10000",x"0C3E2",x"10004",x"0C403",x"10001",x"0C3E3",
									 x"10004",x"0C3E2",x"10008",x"0C3E3",x"10004",x"0C3E2",x"1000A",x"0C3E3",x"10005",x"0CBE3",
									 x"10003",x"0CBE2",x"10004",x"0CC02",x"0C403",x"10002",x"0C3E2",x"10003",x"0BBE2",x"0BBC2",
									 x"10001",x"0B3A2",x"10000",x"0B382",x"0AB61",x"0A342",x"0A322",x"092E2",x"08AE1",x"0A3E2",
									 x"0BD03",x"0DE66",x"0F787",x"0FF87",x"0FF46",x"0FF05",x"0FEE5",x"0FEC5",x"10000",x"0FEA5",
									 x"0FEC5",x"10002",x"0FEA5",x"10001",x"0FE85",x"10002",x"0FE65",x"0FE45",x"10000",x"0FE25",
									 x"0FE24",x"0FE04",x"10000",x"0FDE4",x"0FDC4",x"0FDA4",x"0FD84",x"0FD64",x"0F544",x"0F523",
									 x"0FD02",x"0FCA2",x"0F482",x"0EC43",x"0E4A7",x"0DD2E",x"0DDB3",x"0D637",x"0D69A",x"0DF1C",
									 x"0EF7D",x"0FFDF",x"0FFFF",x"10017",x"0FFFF",x"10018",x"0FFDF",x"0F7DF",x"0EF5D",x"0DEBA",
									 x"0D679",x"0D616",x"0DDB2",x"0DD0C",x"0EC87",x"0EC64",x"0F482",x"0FCC3",x"0F4E4",x"0F524",
									 x"0FD44",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",x"10000",x"0FE04",x"0FE05",x"0FE25",x"0FE45",
									 x"10000",x"0FE65",x"10001",x"0FE85",x"10002",x"0FEA5",x"10002",x"0FEC5",x"10002",x"0FEE5",
									 x"0FF05",x"0FF66",x"0FF87",x"0F767",x"0DE65",x"0B503",x"0AC02",x"09321",x"092E1",x"0A322",
									 x"0AB42",x"0B383",x"0B382",x"10000",x"0B3A2",x"0BBC2",x"10000",x"0BBE2",x"0C3E2",x"10002",
									 x"0C3E3",x"10000",x"0C403",x"0CC03",x"0CC02",x"0C402",x"0CC03",x"10000",x"0C403",x"10000",
									 x"0C3E3",x"0C403",x"10023",x"0C3E2",x"10001",x"0C3E3",x"10001",x"0C403",x"10005",x"0CC03",
									 x"10004",x"0CC02",x"10003",x"0C402",x"0C403",x"10002",x"0C3E2",x"10002",x"0BBE2",x"0BBC2",
									 x"10001",x"0B3A2",x"10000",x"0B382",x"0AB62",x"0A342",x"0A322",x"09B02",x"09301",x"09BA1",
									 x"0C544",x"0DE66",x"0F747",x"0FF86",x"0FF46",x"0FF25",x"0FF05",x"0FEE5",x"0FEC5",x"10000",
									 x"0FEA5",x"0FEC5",x"10002",x"0FEA5",x"10000",x"0FE85",x"10000",x"0FE65",x"10001",x"0FE45",
									 x"10001",x"0FE25",x"0FE04",x"10000",x"0FDE4",x"0FDC4",x"10000",x"0FD84",x"10000",x"0F544",
									 x"0F524",x"0F503",x"0FCC2",x"0FC82",x"0F463",x"0EC66",x"0DCEC",x"0DDD3",x"0D617",x"0CE59",
									 x"0DEDB",x"0EF5D",x"0F7BE",x"0FFDF",x"0FFFF",x"10017",x"0FFFF",x"1001A",x"0F7BF",x"0E71C",
									 x"0D6BA",x"0CE79",x"0D616",x"0D571",x"0E4EB",x"0E486",x"0EC82",x"0F4A2",x"0F4C2",x"0F503",
									 x"0FD44",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"10000",x"0FDE4",x"0FE05",x"0FE25",x"10000",
									 x"0FE45",x"10000",x"0FE65",x"10000",x"0FE85",x"10001",x"0FEA5",x"10002",x"0FEC5",x"10002",
									 x"0FEA5",x"0FEC5",x"0FEE5",x"0FF45",x"0FF66",x"0FFA7",x"0F767",x"0E6C6",x"0CDA5",x"0A3E2",
									 x"09300",x"092E1",x"09B02",x"0AB43",x"0AB42",x"0B382",x"10000",x"0B3A2",x"0BBC2",x"10000",
									 x"0BBE2",x"0C3E2",x"10001",x"0C3E3",x"0C403",x"10000",x"0C402",x"10002",x"0C403",x"0C402",
									 x"0C403",x"10010",x"0CC03",x"10000",x"0C403",x"10001",x"0CC03",x"0C403",x"1001A",x"0CC03",
									 x"10004",x"0CC02",x"10000",x"0C402",x"10000",x"0CC02",x"0C403",x"10001",x"0C3E2",x"10003",
									 x"0BBE2",x"0BBC2",x"10001",x"0B3A2",x"10000",x"0B382",x"0AB62",x"0A342",x"0A322",x"09B02",
									 x"09322",x"09BA1",x"0C544",x"0E6A6",x"0FF88",x"0FF86",x"0FF65",x"0FF05",x"0FEE5",x"10000",
									 x"0FEC5",x"10001",x"0FEA5",x"0FEC5",x"10002",x"0FEA5",x"10000",x"0FE85",x"10000",x"0FE65",
									 x"10001",x"0FE45",x"10000",x"0FE25",x"0FE05",x"0FE04",x"0FDE4",x"10000",x"0FDC4",x"0FDA4",
									 x"0FD84",x"0F564",x"0F543",x"0F504",x"0F4E3",x"0FCA3",x"0F463",x"0F485",x"0E4CA",x"0D570",
									 x"0CE36",x"0CE59",x"0CE9A",x"0E73C",x"0F7BE",x"0FFDF",x"0FFFF",x"10018",x"0FFFF",x"1001A",
									 x"0FFDF",x"0EF7D",x"0DEFB",x"0CE9A",x"0CE37",x"0D5D4",x"0D54F",x"0DCE9",x"0E484",x"0F482",
									 x"0F4A2",x"0F4E3",x"0FD23",x"0FD44",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"10000",x"0FDE5",
									 x"0FE05",x"0FE25",x"0FE45",x"10000",x"0FE65",x"10001",x"0FE85",x"10000",x"0FEA5",x"10002",
									 x"0FEC5",x"10001",x"0FEA5",x"10000",x"0FEC5",x"0FEE5",x"0FF05",x"0FF25",x"0FF66",x"0FF86",
									 x"0F767",x"0E6C6",x"0C544",x"0A3E1",x"09321",x"092C1",x"0A322",x"0AB42",x"0AB62",x"0B382",
									 x"0B3A2",x"0B3C2",x"0BBC2",x"10000",x"0BBE2",x"0C3E2",x"10000",x"0C403",x"10000",x"0C402",
									 x"10001",x"0C403",x"10001",x"0C422",x"10002",x"0C403",x"0CC23",x"10003",x"0C403",x"1000A",
									 x"0C402",x"0CC22",x"10003",x"0CC23",x"10011",x"0C403",x"10004",x"0C402",x"10000",x"0C403",
									 x"10002",x"0C402",x"10003",x"0C403",x"10001",x"0C402",x"10000",x"0C3E2",x"10001",x"0BBE2",
									 x"0BBC2",x"10000",x"0B3C2",x"0B3A2",x"0B382",x"0AB62",x"0A342",x"09B22",x"092E1",x"09301",
									 x"09BE2",x"0B4C2",x"0DE85",x"0F746",x"0FF87",x"0FF46",x"0FF25",x"0FF05",x"0FEE5",x"10000",
									 x"0FEC5",x"10001",x"0FEA5",x"0FEC5",x"10001",x"0FEA5",x"10000",x"0FE85",x"10000",x"0FE65",
									 x"10001",x"0FE45",x"10000",x"0FE25",x"10000",x"0FE05",x"0FDE4",x"10000",x"0FDC4",x"0FDA4",
									 x"10000",x"0FD64",x"0F544",x"0F503",x"0F4E3",x"0F4A3",x"0F463",x"0EC45",x"0E4A8",x"0DD2E",
									 x"0CDD3",x"0CE58",x"0CE99",x"0DEFA",x"0EF9C",x"0FFFF",x"1001A",x"0FFFF",x"1001B",x"0FFBE",
									 x"0E73C",x"0D6BB",x"0CE59",x"0CDF7",x"0CDB3",x"0DD2D",x"0E486",x"0F464",x"0F463",x"0F4A4",
									 x"0FD03",x"0FD23",x"0FD44",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FE05",x"10001",x"0FE25",
									 x"0FE45",x"10000",x"0FE65",x"10000",x"0FE85",x"10000",x"0FEA5",x"10002",x"0FEC5",x"10004",
									 x"0FEE5",x"10001",x"0FF26",x"0FF66",x"0FFA6",x"0F766",x"0E686",x"0BCE3",x"09BC2",x"09301",
									 x"092E1",x"09B22",x"0AB62",x"0ABA2",x"10000",x"0B3A2",x"0B3C2",x"0BBC2",x"0BBE3",x"10000",
									 x"0C3E2",x"10000",x"0C402",x"0C3E2",x"10000",x"0C402",x"10000",x"0C403",x"10000",x"0C423",
									 x"0C422",x"10001",x"0CC22",x"10000",x"0CC23",x"1000E",x"0CC22",x"10004",x"0CC23",x"10016",
									 x"0C402",x"1000A",x"0C403",x"10001",x"0C402",x"10000",x"0C3E2",x"10000",x"0BBE3",x"0BBE2",
									 x"0BBC2",x"0B3C2",x"0B3A2",x"0B382",x"0AB62",x"0A342",x"0A322",x"09B01",x"09301",x"09BA2",
									 x"0B4E4",x"0D625",x"0F786",x"0FF85",x"0FF66",x"0FF26",x"0FF05",x"0FEE5",x"0FEC5",x"0FEC6",
									 x"10000",x"0FEC5",x"10000",x"0FEA5",x"10000",x"0FEC5",x"0FEA5",x"10001",x"0FE85",x"10000",
									 x"0FE65",x"10000",x"0FE45",x"10000",x"0FE25",x"10000",x"0FE05",x"10000",x"0FDE4",x"0FDC4",
									 x"0FDA4",x"0FD84",x"10000",x"0FD44",x"0F523",x"0FCE3",x"0F4C3",x"0F484",x"0F444",x"0E487",
									 x"0DCEB",x"0D592",x"0CE16",x"0CE59",x"0D69A",x"0E71B",x"0EFBE",x"0FFFF",x"1001A",x"0FFFF",
									 x"1001B",x"0FFDF",x"0EF7D",x"0E71C",x"0DEBA",x"0D659",x"0CDF7",x"0D593",x"0DCEC",x"0EC86",
									 x"0F464",x"0F484",x"0FCC3",x"0FD03",x"0FD23",x"0F564",x"0F584",x"0FD84",x"0FDA4",x"0FDE5",
									 x"10000",x"0FE04",x"0FE05",x"0FE25",x"0FE45",x"10000",x"0FE65",x"0FE85",x"10001",x"0FEA5",
									 x"10002",x"0FEC5",x"10002",x"0FEE5",x"10002",x"0FF06",x"0FF26",x"0FF66",x"0FF86",x"0FF87",
									 x"0E6C6",x"0CDA5",x"0AC43",x"09321",x"092C1",x"09AE2",x"0A322",x"0AB62",x"0AB82",x"0B3A2",
									 x"10000",x"0BBA2",x"0BBC2",x"10000",x"0BBE2",x"10001",x"0C402",x"10001",x"0C423",x"10000",
									 x"0C422",x"0CC22",x"10002",x"0CC23",x"10009",x"0C423",x"10000",x"0CC23",x"10002",x"0CC22",
									 x"0CC23",x"10010",x"0C423",x"10000",x"0CC23",x"10007",x"0CC22",x"10001",x"0C423",x"10000",
									 x"0C403",x"0C423",x"0C402",x"10001",x"0C422",x"10000",x"0C423",x"0C403",x"10001",x"0C402",
									 x"0BBE2",x"10000",x"0BBC3",x"0B3C2",x"10000",x"0B3A2",x"0B382",x"0AB62",x"0AB43",x"09AE2",
									 x"092E1",x"09341",x"0AC03",x"0CD85",x"0E6C7",x"0F767",x"0FFA6",x"0FF45",x"0FF25",x"0FF05",
									 x"0FEE5",x"10000",x"0FEC5",x"10004",x"0FEA5",x"10002",x"0FE85",x"10000",x"0FE65",x"10000",
									 x"0FE45",x"10000",x"0FE25",x"10000",x"0FE05",x"10000",x"0FDE5",x"0FDE4",x"0FDA4",x"0FD84",
									 x"0F584",x"0FD64",x"0FD44",x"0FD03",x"0FCC3",x"0FC83",x"0F464",x"0EC46",x"0E4EB",x"0D591",
									 x"0CDF6",x"0CE58",x"0D6BA",x"0E71C",x"0F77D",x"0FFDF",x"0FFFF",x"1001A",x"0FFFF",x"1001C",
									 x"0FFDF",x"0EF7D",x"0E71C",x"0D699",x"0CE38",x"0D5F7",x"0D551",x"0DCC9",x"0EC85",x"0F464",
									 x"0FCA2",x"0FCC2",x"0FD03",x"0F544",x"0F564",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",x"10000",
									 x"0FE04",x"10000",x"0FE25",x"0FE45",x"10000",x"0FE65",x"0FE85",x"10002",x"0FEA5",x"10001",
									 x"0FEC5",x"10002",x"0FEE5",x"10001",x"0FF05",x"0FF25",x"0FF26",x"0FF46",x"0FFA7",x"0F786",
									 x"0E6C5",x"0D5C4",x"0B463",x"09B42",x"09B02",x"10000",x"0A362",x"0AB62",x"0AB82",x"0B382",
									 x"0B3A2",x"0B3C2",x"0BBE2",x"10000",x"0BC02",x"10000",x"0C402",x"0C403",x"0C423",x"0C422",
									 x"0C423",x"0C422",x"0CC23",x"0CC22",x"0C422",x"10000",x"0CC23",x"10008",x"0C423",x"10005",
									 x"0CC23",x"10010",x"0C423",x"10004",x"0CC23",x"10004",x"0CC22",x"10000",x"0CC23",x"10000",
									 x"0C423",x"10001",x"0C422",x"10003",x"0C423",x"0C403",x"0BC02",x"10000",x"0BBE2",x"10001",
									 x"0B3C3",x"0B3C2",x"0ABA2",x"0B3A2",x"0B362",x"0A342",x"09B22",x"09B02",x"09B82",x"0B463",
									 x"0CD85",x"0EEC7",x"0EF67",x"0FF87",x"0FF66",x"0FF25",x"0FF05",x"0FEE5",x"10001",x"0FEC5",
									 x"10004",x"0FEA5",x"10002",x"0FE85",x"10000",x"0FE65",x"10000",x"0FE45",x"0FE25",x"10000",
									 x"0FE05",x"10000",x"0FDE4",x"0FDC4",x"10000",x"0FDA3",x"0FD83",x"0F564",x"0F544",x"0FD03",
									 x"0F4C2",x"0FC82",x"0F463",x"0EC65",x"0E488",x"0DD4F",x"0CDF6",x"0C638",x"0CE79",x"0DEFB",
									 x"0EF5D",x"0F7BE",x"0FFFF",x"1001B",x"0FFFF",x"1001D",x"0F7BE",x"0EF5D",x"0DEDA",x"0CE59",
									 x"0CE58",x"0CDD4",x"0D54E",x"0E4E8",x"0EC85",x"0F483",x"0FCA2",x"0FCC2",x"0F504",x"0F544",
									 x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",x"10000",x"0FE04",x"0FE24",x"0FE25",x"0FE45",
									 x"10000",x"0FE65",x"10000",x"0FE85",x"10001",x"0FEA5",x"10001",x"0FEC5",x"10002",x"0FEE5",
									 x"10000",x"0FF05",x"0FEE5",x"0FF05",x"0FF25",x"0FF66",x"0FFA6",x"0FF87",x"0F747",x"0CDE4",
									 x"0B482",x"09BA1",x"09321",x"09301",x"09B41",x"0AB62",x"0AB82",x"0B3A2",x"0B3C2",x"0B3E2",
									 x"0BBE2",x"10000",x"0BC02",x"10000",x"0C402",x"0C403",x"10000",x"0C423",x"10000",x"0C422",
									 x"10002",x"0CC23",x"10003",x"0CC43",x"10000",x"0CC23",x"10002",x"0CC43",x"1001C",x"0CC23",
									 x"0CC22",x"10004",x"0CC23",x"10003",x"0C423",x"0C403",x"0C423",x"10000",x"0C422",x"10000",
									 x"0C423",x"0BC02",x"10000",x"0BBE2",x"10000",x"0BBC2",x"0B3C2",x"0B3E2",x"0B3C2",x"0AB82",
									 x"0A362",x"0A321",x"09B01",x"09301",x"09BA1",x"0B481",x"0CDA4",x"0EEC6",x"0FF88",x"0FF87",
									 x"0FF66",x"0FF46",x"0FF05",x"0FEE5",x"0FEC5",x"0FEE5",x"10001",x"0FEC5",x"10002",x"0FEA5",
									 x"10002",x"0FE85",x"10000",x"0FE65",x"10000",x"0FE45",x"10000",x"0FE25",x"0FE04",x"10000",
									 x"0FDE4",x"0FDC4",x"10000",x"0FDA4",x"0FD83",x"0FD63",x"0FD43",x"0FD23",x"0FCE3",x"0F482",
									 x"0F483",x"0E485",x"0DCC8",x"0DD2D",x"0D5B3",x"0C658",x"0C679",x"0D6BA",x"0EF5D",x"0F79E",
									 x"0FFDF",x"0FFFF",x"1001B",x"0FFFF",x"1001E",x"0F7BE",x"0E73C",x"0DEBA",x"0CE79",x"0C637",
									 x"0D5D3",x"0DD2E",x"0E4A9",x"0EC85",x"0F483",x"0FCA2",x"0F4E3",x"0F524",x"0FD44",x"0FD64",
									 x"0FDA4",x"10000",x"0FDC4",x"0FDE4",x"10000",x"0FE04",x"10000",x"0FE25",x"0FE45",x"10000",
									 x"0FE65",x"10000",x"0FE85",x"10001",x"0FEA5",x"10000",x"0FEC5",x"10003",x"0FEE5",x"10000",
									 x"0FEC5",x"0FEE5",x"0FF05",x"0FF25",x"0FF45",x"0FFA6",x"0FFE7",x"0F746",x"0DE65",x"0C544",
									 x"0A422",x"09341",x"09301",x"09B02",x"0A343",x"0AB83",x"0ABA2",x"0B3C2",x"10000",x"0B3E2",
									 x"0BBE2",x"10000",x"0BC02",x"10000",x"0C403",x"0C423",x"10000",x"0C422",x"10002",x"0C423",
									 x"10002",x"0CC23",x"0CC43",x"10023",x"0CC22",x"10003",x"0CC42",x"0C443",x"0C423",x"10005",
									 x"0C403",x"0C422",x"10000",x"0BC03",x"0BC02",x"0BBE2",x"10000",x"0BBC2",x"0B3C2",x"10000",
									 x"0ABA2",x"0AB82",x"0A342",x"09B22",x"09301",x"09B62",x"0A3E2",x"0C564",x"0E665",x"0F746",
									 x"0FF87",x"0FFA7",x"0FF66",x"0FF26",x"0FF05",x"0FEE5",x"0FEC5",x"10005",x"0FEA5",x"10003",
									 x"0FE85",x"10000",x"0FE65",x"10000",x"0FE45",x"0FE25",x"10001",x"0FE04",x"0FDE4",x"10000",
									 x"0FDC4",x"0FDA4",x"0FD84",x"0FD64",x"0FD23",x"10000",x"0FCE3",x"0FCA3",x"0F463",x"0EC85",
									 x"0E4A8",x"0DD2D",x"0DDB2",x"0CDF6",x"0C67A",x"0D6BB",x"0E73C",x"0F7BE",x"0FFFF",x"1001D",
									 x"0FFFF",x"1001F",x"0F79E",x"0EEFC",x"0D69A",x"0CE58",x"0D617",x"0DD92",x"0DD0E",x"0E4A8",
									 x"0EC65",x"0FCA3",x"0F4C3",x"0F4E3",x"0FD03",x"0FD44",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",
									 x"0FDE4",x"10000",x"0FE04",x"0FE25",x"0FE45",x"10000",x"0FE65",x"10001",x"0FE85",x"10000",
									 x"0FEA5",x"10001",x"0FEC5",x"10006",x"0FEE5",x"0FF05",x"0FF25",x"0FF86",x"0FFC6",x"10000",
									 x"0FF86",x"0EEC6",x"0CDA5",x"0AC43",x"09B82",x"09322",x"09B22",x"0A343",x"0A363",x"0ABA2",
									 x"0B3A2",x"0B3C2",x"0BBE2",x"10001",x"0BC02",x"0C403",x"0C423",x"0C403",x"10000",x"0C423",
									 x"0C422",x"10000",x"0C423",x"0C422",x"10000",x"0C423",x"10000",x"0CC43",x"10022",x"0CC42",
									 x"0C442",x"10004",x"0C443",x"0C423",x"10000",x"0C443",x"0C423",x"10001",x"0C403",x"0C402",
									 x"0C403",x"0BC02",x"10000",x"0BBE2",x"10000",x"0B3C2",x"10000",x"0B3A2",x"0AB82",x"0A363",
									 x"09B22",x"10000",x"09321",x"09B82",x"0B463",x"0C564",x"0EEC6",x"0F786",x"0FFC6",x"0FFA6",
									 x"0FF45",x"0FF25",x"0FF05",x"0FF06",x"0FEE6",x"0FEC5",x"10004",x"0FEA5",x"10003",x"0FE85",
									 x"10000",x"0FE65",x"10000",x"0FE45",x"0FE25",x"10001",x"0FE05",x"0FDE4",x"0FDC4",x"10000",
									 x"0FDA4",x"0FD84",x"0FD64",x"0FD44",x"0F503",x"0FCE2",x"0FCC3",x"0F483",x"0F464",x"0EC87",
									 x"0DD0C",x"0D592",x"0D616",x"0CE38",x"0D69A",x"0DF1C",x"0EF7D",x"0FFDF",x"0FFFF",x"1001D",
									 x"0FFFF",x"1001F",x"0F7BF",x"0EF5D",x"0DEFA",x"0CE98",x"0CE18",x"0CDD6",x"0D592",x"0DCEC",
									 x"0E487",x"0F484",x"0F4A3",x"0F4C3",x"0F4E3",x"0F523",x"0FD44",x"0FD64",x"0FD84",x"0FDA4",
									 x"0FDC4",x"0FDE4",x"10000",x"0FE05",x"0FE25",x"10000",x"0FE45",x"10000",x"0FE65",x"0FE85",
									 x"10002",x"0FEA5",x"10000",x"0FEC5",x"10002",x"0FEE5",x"10003",x"0FF06",x"0FF26",x"0FF46",
									 x"0FFA6",x"0FFA7",x"0F767",x"0EEE6",x"0CDC4",x"0BCC4",x"0AC02",x"09301",x"092E1",x"09B22",
									 x"0A362",x"0ABA2",x"10000",x"0B3C2",x"0B3E2",x"0BBE2",x"0BC02",x"0BC03",x"10000",x"0BC02",
									 x"0C402",x"10000",x"0C422",x"10000",x"0C423",x"0C422",x"10000",x"0C423",x"10000",x"0CC43",
									 x"10022",x"0CC42",x"0C442",x"10004",x"0C443",x"0C423",x"10003",x"0C403",x"10000",x"0BC02",
									 x"0BC03",x"0BC02",x"10001",x"0B3E2",x"0B3C2",x"0ABA2",x"0AB82",x"0A362",x"09B21",x"09301",
									 x"09B41",x"0A3C1",x"0BCE4",x"0D5E5",x"0E6E5",x"0F767",x"0FFA6",x"10000",x"0FF26",x"0FF05",
									 x"10000",x"0FEE5",x"0FEE6",x"10000",x"0FEE5",x"0FEC5",x"10002",x"0FEA5",x"10003",x"0FE85",
									 x"10001",x"0FE65",x"0FE45",x"10000",x"0FE25",x"10000",x"0FE05",x"0FDE5",x"0FDC4",x"10000",
									 x"0FDA4",x"0FD84",x"0FD63",x"0FD43",x"0FD24",x"0FCE3",x"0FCC2",x"0F4A3",x"0EC64",x"0EC66",
									 x"0E4CA",x"0DD90",x"0CE16",x"0C638",x"0CE79",x"0DEFB",x"0EF5C",x"0F7BE",x"0FFFF",x"1001E",
									 x"0FFFF",x"10020",x"0F7BE",x"0EF7C",x"0DEFA",x"0CE79",x"0CE38",x"0CDF5",x"0D570",x"0DCEB",
									 x"0EC86",x"0F464",x"0F4A3",x"0F4C3",x"0F503",x"0F543",x"0F563",x"0F584",x"0FD84",x"0FDA4",
									 x"0FDC4",x"10000",x"0FDE5",x"0FE05",x"0FE25",x"10000",x"0FE45",x"0FE65",x"0FE85",x"10002",
									 x"0FEA5",x"10001",x"0FEC5",x"10001",x"0FEE5",x"10000",x"0FEE6",x"10001",x"0FF06",x"10000",
									 x"0FF26",x"0FF66",x"0FF86",x"0FF87",x"0FFA7",x"0EF06",x"0DE45",x"0C563",x"0AC41",x"09B81",
									 x"09B42",x"09301",x"09B41",x"0A361",x"0B3A2",x"0B3C2",x"0B3E2",x"10000",x"0BBE3",x"0BC02",
									 x"10002",x"0C422",x"0C423",x"10004",x"0C443",x"0CC43",x"10007",x"0C443",x"0CC43",x"10017",
									 x"0CC42",x"0C442",x"10003",x"0C443",x"10000",x"0C423",x"10002",x"0C403",x"0BC03",x"0BC02",
									 x"10001",x"0B402",x"0B3E2",x"0B3C2",x"10000",x"0B3C3",x"0A362",x"09B01",x"10000",x"09321",
									 x"09BA1",x"0AC41",x"0BD23",x"0DE66",x"0F727",x"0FFA7",x"0FFC7",x"0FF86",x"0FF46",x"0FF06",
									 x"0FEE5",x"10001",x"0FEE6",x"10000",x"0FEE5",x"0FEC5",x"10001",x"0FEA5",x"10002",x"0FE85",
									 x"10001",x"0FE65",x"10001",x"0FE45",x"0FE25",x"10000",x"0FE05",x"10000",x"0FDE4",x"0FDC4",
									 x"0FDA4",x"0FD84",x"10000",x"0FD44",x"0FD23",x"0FD03",x"0FCC2",x"0F4A2",x"0F483",x"0E486",
									 x"0E4CA",x"0D54E",x"0CDD4",x"0C637",x"0C699",x"0D6FA",x"0EF5C",x"0F79E",x"0FFDF",x"0FFFF",
									 x"1001E",x"0FFFF",x"10021",x"0F7BE",x"0EF5C",x"0DEFA",x"0CE79",x"0CE38",x"0CDD4",x"0D571",
									 x"0ECEB",x"0F487",x"0F464",x"0F483",x"0F4C2",x"0F502",x"0F543",x"0F544",x"0F564",x"0FD83",
									 x"0FDA4",x"0FDC4",x"0FDC5",x"0FDE5",x"0FE05",x"0FE25",x"10000",x"0FE45",x"0FE65",x"0FE85",
									 x"10003",x"0FEA5",x"10000",x"0FEC5",x"10002",x"0FEE5",x"10003",x"0FF05",x"0FF26",x"0FF46",
									 x"0FF45",x"0FF86",x"0FFA6",x"0FFA7",x"0F746",x"0D665",x"0C544",x"0B443",x"0A382",x"09321",
									 x"09B41",x"0A341",x"0AB62",x"0ABA2",x"10000",x"0B3C2",x"0B3E2",x"0B402",x"0BC02",x"0BC03",
									 x"10000",x"0BC22",x"0BC23",x"0C423",x"10004",x"0C442",x"10001",x"0C443",x"10006",x"0CC43",
									 x"10010",x"0C443",x"10007",x"0C442",x"0C422",x"0C443",x"10000",x"0C423",x"10002",x"0BC03",
									 x"10000",x"0BC02",x"0B402",x"0B3E2",x"10000",x"0B3C2",x"0ABA2",x"0AB82",x"0A362",x"09B21",
									 x"09321",x"09B41",x"0AC22",x"0C564",x"0D645",x"0EF26",x"0FFA8",x"0FFA7",x"10000",x"0FF66",
									 x"0FF25",x"0FF05",x"0FEE5",x"10000",x"0FEC5",x"0FEE5",x"10000",x"0FEC5",x"10002",x"0FEA5",
									 x"10001",x"0FE85",x"10002",x"0FE65",x"10001",x"0FE45",x"0FE25",x"10000",x"0FE04",x"0FE05",
									 x"0FDE4",x"0FDC4",x"0FDA4",x"0FD84",x"10000",x"0FD64",x"0FD23",x"0FCE3",x"0FCC3",x"0FC82",
									 x"0F462",x"0EC85",x"0E4EB",x"0D570",x"0CDD4",x"0D637",x"0D679",x"0D6DA",x"0E75C",x"0F7BE",
									 x"0FFDF",x"0FFFF",x"1001F",x"0FFFF",x"10022",x"0F7BE",x"0E73C",x"0D6BA",x"0CE79",x"0C5F7",
									 x"0CDB4",x"0DD51",x"0E4CB",x"0EC66",x"0F464",x"0F483",x"0F4C2",x"0FD02",x"0F523",x"0F564",
									 x"0FD83",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",x"0FE04",x"10000",x"0FE24",x"0FE45",x"0FE65",
									 x"10001",x"0FE85",x"10002",x"0FEA5",x"10000",x"0FEC5",x"10003",x"0FEE5",x"10001",x"0FF05",
									 x"10000",x"0FF25",x"0FF46",x"10000",x"0FF65",x"0FFA6",x"0FFC6",x"0F786",x"0E6E6",x"0DE25",
									 x"0C544",x"0AC22",x"09B82",x"09301",x"09B02",x"0A362",x"0AB82",x"0ABA1",x"0B3C2",x"10000",
									 x"0B3C3",x"0BBE4",x"0BBE3",x"0BC02",x"10000",x"0BC22",x"10000",x"0C422",x"10000",x"0C423",
									 x"10000",x"0C443",x"0C442",x"10000",x"0C443",x"10006",x"0CC43",x"1000F",x"0C443",x"1000A",
									 x"0C422",x"10000",x"0BC22",x"10000",x"0BC23",x"0BC02",x"10000",x"0B402",x"0B3E3",x"0B3C3",
									 x"10000",x"0B3A3",x"0A361",x"09B21",x"09301",x"08B00",x"09BA1",x"0AC62",x"0C523",x"0D605",
									 x"0EF07",x"0F766",x"0FFA6",x"0FF86",x"0FF66",x"0FF46",x"0FF26",x"0FF05",x"0FEE5",x"0FEC5",
									 x"10005",x"0FEA5",x"10002",x"0FE85",x"10001",x"0FE65",x"10001",x"0FE45",x"10000",x"0FE25",
									 x"10000",x"0FE04",x"0FDE4",x"10000",x"0FDC4",x"0FDA4",x"0FD84",x"0F584",x"0F543",x"0F523",
									 x"0FD03",x"0FCC2",x"0F483",x"0F463",x"0EC65",x"0E4CA",x"0D54F",x"0CDB4",x"0CDF6",x"0CE59",
									 x"0D6BB",x"0E73C",x"0F79D",x"0FFDE",x"0FFFF",x"10020",x"0FFFF",x"10022",x"0FFDE",x"0EF9D",
									 x"0E73C",x"0D6BA",x"0C638",x"0C5F7",x"0CDB4",x"0D52F",x"0E4A9",x"0EC65",x"0F464",x"0F4A3",
									 x"0FCC2",x"0FCE3",x"0F523",x"0F564",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",x"0FE04",
									 x"0FE05",x"0FE25",x"0FE45",x"0FE65",x"10002",x"0FE85",x"10001",x"0FEA5",x"10001",x"0FEC5",
									 x"10002",x"0FEE5",x"0FEC5",x"0FEE5",x"10001",x"0FF05",x"0FF25",x"0FF46",x"0FF86",x"0FFC7",
									 x"0FFE7",x"0FFA7",x"0EF26",x"0DE64",x"0C583",x"0AC83",x"09BA2",x"09322",x"09B21",x"09B42",
									 x"0A362",x"0AB82",x"0ABA3",x"0B3A2",x"0B3C3",x"0B3E3",x"0B3E2",x"0BC02",x"10000",x"0BC22",
									 x"10001",x"0BC23",x"0C423",x"0C443",x"1000A",x"0CC43",x"1000A",x"0C443",x"0CC43",x"10001",
									 x"0C443",x"10009",x"0C423",x"0BC22",x"10001",x"0BC02",x"0BC03",x"10000",x"0B402",x"0B3E2",
									 x"0B3C3",x"0ABA3",x"0AB82",x"0AB62",x"0A342",x"09B22",x"09301",x"09361",x"0AC42",x"0C563",
									 x"0DE65",x"0EF06",x"0FFA7",x"10000",x"0FFA6",x"0FF66",x"0FF45",x"0FF26",x"0FEE5",x"10002",
									 x"0FEC5",x"10002",x"0FEA5",x"10003",x"0FE85",x"10001",x"0FE65",x"10002",x"0FE45",x"0FE25",
									 x"10000",x"0FE05",x"0FDE4",x"10000",x"0FDC4",x"0FDA4",x"0FD84",x"10000",x"0F564",x"0F523",
									 x"0F502",x"0FCC2",x"0F4A2",x"0F483",x"0EC85",x"0E4C9",x"0D52E",x"0CDB3",x"0C5F6",x"0C637",
									 x"0D69A",x"0E71D",x"0EF7D",x"0FFDE",x"0FFDF",x"0FFFF",x"10020",x"0FFFF",x"10023",x"0FFDE",
									 x"0F79E",x"0E71C",x"0CEBA",x"0C658",x"0C616",x"0CDB3",x"0DD4E",x"0DCCA",x"0E487",x"0EC84",
									 x"0FCA3",x"10000",x"0FCE3",x"0F524",x"0FD44",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",
									 x"0FE04",x"0FE05",x"0FE25",x"0FE45",x"10000",x"0FE65",x"10002",x"0FE85",x"10000",x"0FEA5",
									 x"10002",x"0FEC5",x"0FEC6",x"10000",x"0FEC5",x"10001",x"0FEE5",x"10000",x"0FF05",x"10000",
									 x"0FF26",x"0FF46",x"0FF86",x"0FF87",x"10000",x"0F767",x"0EF07",x"0DE66",x"0CD85",x"0B483",
									 x"09BA0",x"09340",x"09321",x"09B42",x"0A382",x"0AB82",x"0ABA2",x"0B3C2",x"0B3E3",x"0B403",
									 x"10000",x"0BC03",x"0BC22",x"10000",x"0BC23",x"10001",x"0BC43",x"10000",x"0C443",x"0C423",
									 x"10002",x"0C443",x"10015",x"0C422",x"0C443",x"0C422",x"0C423",x"0C443",x"0C423",x"10000",
									 x"0BC23",x"10000",x"0BC22",x"10000",x"0B402",x"0B403",x"0B3E3",x"0B3C3",x"0ABC2",x"0ABA2",
									 x"0A382",x"0A362",x"09B21",x"09300",x"09320",x"0A3C2",x"0B444",x"0C525",x"0DE47",x"0EF07",
									 x"0F787",x"0FF87",x"0FFA7",x"0FF66",x"0FF46",x"0FF06",x"0FF05",x"10000",x"0FEE5",x"0FEC5",
									 x"10004",x"0FEA5",x"10003",x"0FE85",x"10001",x"0FE65",x"10001",x"0FE45",x"10000",x"0FE25",
									 x"10000",x"0FE05",x"0FDE5",x"0FDE4",x"0FDC4",x"0FDA4",x"10000",x"0FD84",x"0FD44",x"0FD23",
									 x"0FD03",x"0FCE3",x"0F4A3",x"0F483",x"0ECA5",x"0E4E9",x"0D54E",x"0CDB3",x"0C616",x"0C658",
									 x"0D699",x"0E71C",x"0EF7E",x"0F7BE",x"0FFFF",x"10022",x"0FFFF",x"10023",x"0FFDF",x"10000",
									 x"0F77E",x"0E71B",x"0D69A",x"0CE38",x"0CDD6",x"0D5B3",x"0D550",x"0DCEB",x"0E486",x"0F484",
									 x"0FC63",x"0FCA3",x"0F4E3",x"0F503",x"0FD23",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",
									 x"0FE04",x"10000",x"0FE25",x"10000",x"0FE45",x"10000",x"0FE65",x"10000",x"0FE85",x"10002",
									 x"0FEA5",x"10001",x"0FEC5",x"10006",x"0FEE5",x"10000",x"0FF05",x"0FF26",x"0FF46",x"0FF86",
									 x"0FFA7",x"0FFC7",x"0FFA7",x"0F747",x"0DE66",x"0CD84",x"0BCE4",x"0B464",x"0A3E2",x"09B62",
									 x"09B42",x"09B21",x"0A342",x"0A362",x"0ABA2",x"0ABC2",x"0B3E2",x"10000",x"0B402",x"0BC03",
									 x"0B402",x"0BC03",x"0BC23",x"10000",x"0BC22",x"10003",x"0BC23",x"0C443",x"10012",x"0C442",
									 x"10000",x"0C422",x"0BC22",x"10000",x"0BC23",x"10000",x"0BC02",x"10002",x"0B3E2",x"10000",
									 x"0B3C2",x"0ABC2",x"0ABA2",x"0A362",x"0A342",x"09B42",x"09321",x"09B62",x"0A3E2",x"0AC42",
									 x"0C504",x"0D5A6",x"0DE46",x"0EEE6",x"0FF87",x"0FFC7",x"10000",x"0FF86",x"0FF66",x"0FF26",
									 x"0FF06",x"0FEE5",x"0FEC5",x"10006",x"0FEA5",x"10003",x"0FE85",x"10001",x"0FE65",x"10000",
									 x"0FE45",x"10000",x"0FE25",x"10001",x"0FE05",x"10000",x"0FDE4",x"0FDC4",x"0FDA4",x"0FD84",
									 x"0FD64",x"0F543",x"0FD04",x"0FCE3",x"0FCC3",x"0F4A3",x"0F484",x"0EC85",x"0E4C9",x"0DD4E",
									 x"0D5B3",x"0C5F7",x"0C638",x"0D699",x"0DEFB",x"0EF7E",x"0FFDF",x"0FFFF",x"10023",x"0FFFF",
									 x"10025",x"0FFDF",x"0EF5D",x"0DEFB",x"0D679",x"0CE18",x"0CDF6",x"0CDB4",x"0DD4E",x"0E4A9",
									 x"0F464",x"0FC43",x"0FC83",x"0FCC3",x"0FD03",x"0FD23",x"0F543",x"0F583",x"0FDA4",x"0FDC4",
									 x"10000",x"0FDE4",x"10000",x"0FE04",x"0FE25",x"10001",x"0FE45",x"0FE65",x"10001",x"0FE85",
									 x"10001",x"0FEA5",x"10003",x"0FEC5",x"10003",x"0FEE5",x"10001",x"0FF05",x"0FF26",x"0FF46",
									 x"0FF66",x"0FFA6",x"0FFC6",x"10000",x"0F766",x"0EF06",x"0E6A6",x"0CDA4",x"0AC62",x"09BA1",
									 x"09341",x"092E2",x"09322",x"09B42",x"0A383",x"0ABA3",x"0ABC3",x"0B3C2",x"10000",x"0B3E2",
									 x"10000",x"0B402",x"10000",x"0B422",x"0BC22",x"0BC02",x"0BC22",x"10001",x"0BC42",x"0BC43",
									 x"0BC23",x"0C443",x"10004",x"0C423",x"10000",x"0C443",x"10002",x"0C423",x"10002",x"0C422",
									 x"10000",x"0BC22",x"10000",x"0C422",x"0BC22",x"10000",x"0BC02",x"0BC03",x"0B402",x"0B3E3",
									 x"0BC03",x"0B3E3",x"0B3C2",x"0B3E3",x"0ABC3",x"0ABA2",x"0A362",x"09B42",x"09B01",x"092E1",
									 x"09300",x"09BC1",x"0B4A3",x"0C564",x"0DE66",x"0F726",x"0FF86",x"0FFC6",x"10000",x"0FFA5",
									 x"0FF86",x"0FF45",x"0FF25",x"0FF05",x"0FEE5",x"0FEC5",x"10002",x"0FEA5",x"10007",x"0FE85",
									 x"10001",x"0FE65",x"10000",x"0FE45",x"10001",x"0FE25",x"10000",x"0FE05",x"10000",x"0FDE4",
									 x"0FDC4",x"10000",x"0FD84",x"10000",x"0F563",x"0F543",x"0FD03",x"0FCC3",x"0F482",x"0F483",
									 x"0EC65",x"0E4A7",x"0D52D",x"0D592",x"0CDF6",x"0C619",x"0CE7A",x"0DEDB",x"0EF5C",x"0FFBE",
									 x"0FFFF",x"10024",x"0FFFF",x"10026",x"0F7BE",x"0EF5C",x"0DEDB",x"0D679",x"0CE17",x"0CDF6",
									 x"0D593",x"0DD0D",x"0E488",x"0EC65",x"0F484",x"0F4A3",x"0FCC3",x"0FD03",x"0F522",x"0F543",
									 x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",x"10000",x"0FE04",x"0FE05",x"0FE25",x"10000",
									 x"0FE45",x"10001",x"0FE65",x"10001",x"0FE85",x"10000",x"0FEA5",x"10002",x"0FEC5",x"10003",
									 x"0FEE5",x"10000",x"0FF05",x"10001",x"0FF26",x"0FF66",x"0FF86",x"0FFA6",x"0FFC6",x"0FFA6",
									 x"0F786",x"0EF06",x"0DE44",x"0CDC4",x"0C524",x"0AC63",x"0A3E2",x"09B82",x"09321",x"092E1",
									 x"09B01",x"0A321",x"0AB82",x"0ABA2",x"0B3C2",x"0B3E2",x"10001",x"0B402",x"0B403",x"10001",
									 x"0BC23",x"10012",x"0BC02",x"0BC03",x"10001",x"0B3E3",x"10000",x"0B3E2",x"0B402",x"0B3E2",
									 x"10000",x"0B3E3",x"0B3C3",x"0ABA2",x"0AB82",x"0A342",x"09B00",x"092E0",x"09320",x"09B61",
									 x"0ABE3",x"0B443",x"0BCE3",x"0CDC4",x"0DE65",x"0E6E6",x"0F786",x"0FFC6",x"10000",x"0FFA6",
									 x"0FF86",x"0FF45",x"0FF25",x"0FF05",x"0FEE5",x"10000",x"0FEC5",x"10004",x"0FEA5",x"10003",
									 x"0FE85",x"10002",x"0FE65",x"10000",x"0FE45",x"10001",x"0FE25",x"10000",x"0FE05",x"10001",
									 x"0FDE4",x"0FDC4",x"0FDA4",x"10000",x"0FD64",x"0FD44",x"0F523",x"0F503",x"0F4E3",x"0F4A3",
									 x"0F463",x"0EC85",x"0E4A8",x"0DD0C",x"0D592",x"0CDF5",x"0CE17",x"0CE59",x"0D6DB",x"0EF5D",
									 x"0F79E",x"0FFDF",x"0FFFF",x"10024",x"0FFFF",x"10027",x"0FFDE",x"0EF7D",x"0DEFC",x"0D69A",
									 x"0CE39",x"0CDF7",x"0CD93",x"0D52E",x"0DCEB",x"0E4A7",x"0EC84",x"0F4A3",x"0F4C2",x"0F502",
									 x"0FD03",x"0FD24",x"0FD44",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FDE4",x"10000",x"0FE05",
									 x"0FE25",x"10000",x"0FE45",x"10001",x"0FE65",x"10001",x"0FE85",x"10001",x"0FEA5",x"10002",
									 x"0FEC5",x"10004",x"0FEE5",x"0FF05",x"10001",x"0FF25",x"0FF45",x"0FF66",x"0FF87",x"0FFA6",
									 x"0FFC7",x"0FFA7",x"0FF67",x"0F707",x"0DE65",x"0CDA4",x"0BD04",x"0A442",x"09BC2",x"09B82",
									 x"0A383",x"0A363",x"0A362",x"10002",x"0AB82",x"10000",x"0ABA3",x"0B3C3",x"10000",x"0B3E3",
									 x"10001",x"0BBE2",x"0BC02",x"10000",x"0BBE2",x"0BC02",x"10006",x"0B402",x"10004",x"0B3E3",
									 x"10000",x"0ABE3",x"0ABC3",x"10000",x"0ABA3",x"0ABA2",x"0AB82",x"0A382",x"0A362",x"10003",
									 x"0A3A2",x"0A3C2",x"0AC42",x"0B4C3",x"0CDC5",x"0DE45",x"0EF06",x"0FF87",x"0FFA7",x"0F7A6",
									 x"0FFA6",x"0FF87",x"0FF86",x"0FF46",x"0FF26",x"0FF05",x"0FEE5",x"10001",x"0FEC5",x"10003",
									 x"0FEA5",x"10005",x"0FE85",x"10001",x"0FE65",x"10000",x"0FE45",x"10000",x"0FE25",x"10000",
									 x"0FE05",x"10001",x"0FDE4",x"10000",x"0FDC4",x"0FDA4",x"0FD84",x"0FD64",x"0F544",x"0F523",
									 x"0FD03",x"0FCC2",x"0F482",x"0F463",x"0EC86",x"0E4CA",x"0D50E",x"0D572",x"0CDD5",x"0CE37",
									 x"0CE79",x"0DEDB",x"0EF5D",x"0F7BE",x"0FFFF",x"10026",x"0FFFF",x"10027",x"0FFDF",x"0F7BE",
									 x"0E75D",x"0DF1C",x"0CE9A",x"0C638",x"0C5D6",x"0CDB3",x"0D590",x"0DCEB",x"0EC66",x"0F464",
									 x"0FC82",x"0FCC2",x"0FCE3",x"0F503",x"0F543",x"0FD63",x"0FD84",x"0FDA4",x"0FDC4",x"10000",
									 x"0FDE4",x"10000",x"0FE04",x"0FE05",x"0FE25",x"10000",x"0FE45",x"10001",x"0FE65",x"10000",
									 x"0FE85",x"10001",x"0FEA5",x"10002",x"0FEC5",x"10005",x"0FEE5",x"10000",x"0FF05",x"10000",
									 x"0FF26",x"0FF46",x"0FF66",x"0FF86",x"0FFA6",x"10001",x"0F785",x"0EF45",x"0EF07",x"0DE66",
									 x"0CDC5",x"0C525",x"0B484",x"0A3C3",x"09B42",x"09301",x"10000",x"09B01",x"09B22",x"0A342",
									 x"0A381",x"0A3A1",x"0A3A2",x"0ABA2",x"0ABC2",x"10000",x"0B3C3",x"10003",x"0B3E3",x"10005",
									 x"0B3C3",x"10004",x"0B3C2",x"0ABC2",x"10000",x"0ABA2",x"0A381",x"10000",x"0A362",x"09B22",
									 x"09301",x"09300",x"10000",x"09B61",x"0A3E2",x"0B463",x"0C525",x"0D5C5",x"0DE46",x"0E6C6",
									 x"0F766",x"0F786",x"0FFC6",x"10001",x"0FFA6",x"0FF66",x"0FF46",x"0FF26",x"0FF06",x"0FEE5",
									 x"0FEC5",x"10000",x"0FEE5",x"0FEC5",x"10004",x"0FEA5",x"10003",x"0FE85",x"10001",x"0FE65",
									 x"10001",x"0FE45",x"10000",x"0FE25",x"10000",x"0FE05",x"0FE04",x"0FDE5",x"0FDE4",x"0FDC4",
									 x"10000",x"0FDA3",x"0FD83",x"0FD64",x"0F543",x"0F523",x"0F503",x"0FCC2",x"0FC82",x"0F462",
									 x"0EC85",x"0E4EA",x"0DD4F",x"0CD93",x"0C5D6",x"0C617",x"0CE79",x"0DEFB",x"0E75D",x"0F7BE",
									 x"0FFDF",x"0FFFF",x"10026",x"0FFFF",x"10027",x"0FFDF",x"10000",x"0EF9E",x"0E75D",x"0DEFC",
									 x"0CE7A",x"0C5F7",x"0C5D6",x"0CDB3",x"0D52E",x"0E4AA",x"0EC46",x"0F464",x"0FCA3",x"0F4C2",
									 x"0F502",x"0F543",x"10000",x"0FD44",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FDE4",x"10000",
									 x"0FE04",x"0FE05",x"0FE25",x"10000",x"0FE45",x"10001",x"0FE65",x"10000",x"0FE85",x"10000",
									 x"0FEA5",x"10003",x"0FEC5",x"10006",x"0FEE5",x"0FEE6",x"0FF06",x"10000",x"0FF26",x"0FF46",
									 x"0FF66",x"0FF86",x"0FFC6",x"10002",x"0F766",x"0E6E5",x"0DE65",x"0CDC4",x"0BD23",x"0B484",
									 x"0AC43",x"0A402",x"0A3C2",x"0A3A2",x"10000",x"09B82",x"09B62",x"10000",x"09B42",x"10001",
									 x"0A362",x"10000",x"0A382",x"0A383",x"10000",x"0AB83",x"10000",x"0ABA3",x"10002",x"0AB83",
									 x"10000",x"0AB82",x"0AB62",x"0A362",x"10000",x"0A342",x"0A322",x"0A342",x"09B42",x"09B41",
									 x"09B62",x"0A382",x"0A3A2",x"0A3C2",x"10000",x"0A3E2",x"0AC42",x"0B4C4",x"0C543",x"0CDC3",
									 x"0DE65",x"0EEE6",x"0F746",x"0F786",x"0FFC6",x"10000",x"0FFA6",x"10000",x"0FF86",x"0FF46",
									 x"0FF26",x"0FF06",x"0FEE6",x"0FEC5",x"10006",x"0FEC6",x"10000",x"0FEA6",x"0FEA5",x"10001",
									 x"0FE85",x"10002",x"0FE65",x"10000",x"0FE45",x"10001",x"0FE25",x"10000",x"0FE05",x"0FDE5",
									 x"10000",x"0FDC4",x"10000",x"0FDA4",x"0FD84",x"10000",x"0FD63",x"0FD43",x"0FD22",x"0F4E2",
									 x"0FCC2",x"0F482",x"0F483",x"0E485",x"0DCC9",x"0D52E",x"0CDB3",x"0C5F5",x"0BE17",x"0C659",
									 x"0D6DB",x"0E75D",x"0EF9E",x"0FFDF",x"0FFFF",x"10027",x"0FFFF",x"10029",x"0FFDF",x"0F7BE",
									 x"0EF7D",x"0E6FC",x"0D659",x"0C617",x"0C5D6",x"0CD93",x"0DD50",x"0E4EC",x"0E4A9",x"0EC85",
									 x"0F463",x"0F4A3",x"0F4E2",x"0F503",x"0F524",x"0FD44",x"0FD64",x"0FD83",x"0FDA3",x"0FDC4",
									 x"10000",x"0FDE4",x"0FE04",x"0FE05",x"10000",x"0FE25",x"0FE45",x"10002",x"0FE65",x"0FE85",
									 x"10002",x"0FEA5",x"10001",x"0FEC5",x"10006",x"0FEC6",x"0FEE6",x"0FEE5",x"0FF05",x"0FF06",
									 x"0FF26",x"10000",x"0FF46",x"0FF66",x"0FFA6",x"0FFC6",x"10001",x"0FFC7",x"0FF87",x"0FF67",
									 x"0F748",x"0EF07",x"0E686",x"0D5E5",x"0CD64",x"0BCE3",x"0AC63",x"0A402",x"09BC2",x"09BA1",
									 x"09B61",x"09341",x"09B41",x"10000",x"09B61",x"10005",x"09B62",x"09B61",x"10001",x"09B60",
									 x"09B40",x"09B60",x"10000",x"09B40",x"09B41",x"10000",x"09B61",x"0A3C1",x"0A402",x"0AC63",
									 x"0BCE3",x"0CD84",x"0D605",x"0DE66",x"0EEE7",x"0F768",x"0FF88",x"0FF87",x"0FFA7",x"0FFC7",
									 x"10000",x"0FFA6",x"0FF86",x"0FF66",x"10000",x"0FF45",x"0FF25",x"0FF06",x"10000",x"0FEE5",
									 x"10000",x"0FEC5",x"10003",x"0FEA5",x"10003",x"0FEA6",x"0FEA5",x"10000",x"0FE85",x"10002",
									 x"0FE65",x"0FE45",x"10000",x"0FE25",x"10001",x"0FE05",x"0FE04",x"0FDE5",x"10000",x"0FDC4",
									 x"0FDA4",x"10000",x"0FD84",x"0FD64",x"0FD44",x"0F524",x"0F523",x"0FCE3",x"0FC83",x"0F463",
									 x"0EC65",x"0E4A7",x"0DCEB",x"0D52F",x"0CDB3",x"0C5D6",x"0C617",x"0CE58",x"0DEDB",x"0E75D",
									 x"0F7BE",x"0FFDF",x"0FFFF",x"10028",x"0FFFF",x"1002A",x"0FFDF",x"0F7BE",x"0EF7D",x"0DEDB",
									 x"0CE79",x"0C638",x"0C5F6",x"0CDB4",x"0D572",x"0DD0D",x"0E488",x"0F466",x"0FC64",x"0FC62",
									 x"0FCC2",x"0FCE3",x"0FD24",x"0F544",x"0FD63",x"0FD83",x"0FDA4",x"10000",x"0FDC4",x"10000",
									 x"0FDE4",x"10000",x"0FE04",x"0FE05",x"0FE25",x"0FE24",x"0FE45",x"10000",x"0FE65",x"10001",
									 x"0FE85",x"10001",x"0FEA5",x"10001",x"0FEC5",x"10004",x"0FEC6",x"0FEC5",x"0FEE5",x"10002",
									 x"0FF05",x"10000",x"0FF25",x"0FF46",x"0FF67",x"0FF86",x"10000",x"0FFA6",x"10000",x"0FFC6",
									 x"0FFC5",x"0FFC6",x"0F786",x"0F746",x"0EF06",x"0E6C6",x"0DE65",x"0DE45",x"0DE25",x"0D5C5",
									 x"0CD84",x"0CD64",x"0CD25",x"0C504",x"0BCC3",x"0BCA3",x"0B483",x"10007",x"0B4A3",x"0B4C3",
									 x"0BCC3",x"0BD04",x"0C524",x"0C564",x"0CD84",x"0CDC5",x"0D605",x"0D645",x"0DE85",x"0E6C6",
									 x"0EF06",x"0F746",x"0F786",x"0F7A6",x"0F7C6",x"0FFC6",x"0FFC7",x"0FFC6",x"0FFA7",x"0FF86",
									 x"0FF66",x"0FF46",x"0FF26",x"0FF25",x"0FEE5",x"10000",x"0FEC5",x"0FEE5",x"10000",x"0FEC5",
									 x"10004",x"0FEA5",x"10002",x"0FE85",x"10003",x"0FE65",x"10001",x"0FE45",x"0FE24",x"10000",
									 x"0FE04",x"10001",x"0FDE4",x"0FDC4",x"10001",x"0FDA4",x"0FD84",x"0FD64",x"10000",x"0FD44",
									 x"0F504",x"0F4E4",x"0F4E3",x"0F483",x"0FC44",x"0F445",x"0E488",x"0DCEC",x"0D551",x"0D594",
									 x"0C5D6",x"0C618",x"0CE59",x"0DEDA",x"0EF5D",x"0F7BE",x"0FFDF",x"0FFFF",x"10029",x"0FFFF",
									 x"1002B",x"0FFDF",x"0F7BE",x"0E75C",x"0DEDA",x"0CE99",x"0C638",x"0BDF7",x"0C5D5",x"0D592",
									 x"0DD0D",x"0E4A9",x"0EC86",x"0FC63",x"0FC82",x"0FCC2",x"0F503",x"0F523",x"0F543",x"0FD43",
									 x"0FD64",x"0FD84",x"0FDA4",x"10000",x"0FDC4",x"0FDE5",x"0FDE4",x"0FE04",x"0FE25",x"10000",
									 x"0FE45",x"10002",x"0FE65",x"10000",x"0FE85",x"10001",x"0FEA5",x"10006",x"0FEC5",x"10001",
									 x"0FEE5",x"10005",x"0FF05",x"0FF26",x"0FF46",x"0FF86",x"10000",x"0FFA6",x"0FFC6",x"10001",
									 x"0FFC7",x"10001",x"0FFA7",x"0FF87",x"0F767",x"10000",x"0EF27",x"0EF06",x"0E6A6",x"0DE65",
									 x"0D625",x"0D604",x"0CDE4",x"0CDC4",x"10000",x"0CDA4",x"10001",x"0CDC4",x"10000",x"0CDC5",
									 x"0CDE5",x"0D605",x"0D625",x"0DE65",x"0E6A6",x"0E706",x"0EF46",x"10000",x"0F787",x"0F7A7",
									 x"0FFA7",x"10001",x"0FFC7",x"10000",x"0FFC6",x"10000",x"0FFA6",x"10000",x"0FF66",x"0FF45",
									 x"0FF25",x"0FF06",x"0FEE5",x"10001",x"0FEC5",x"10005",x"0FEA5",x"10000",x"0FEC5",x"0FEA5",
									 x"10001",x"0FE85",x"10002",x"0FE65",x"10003",x"0FE45",x"10000",x"0FE25",x"0FE05",x"0FE04",
									 x"10000",x"0FDE4",x"0FDC4",x"10001",x"0FDA4",x"0FD84",x"0FD64",x"0FD44",x"0FD43",x"0FD23",
									 x"0F4E4",x"0F4C3",x"0F4A2",x"0F463",x"0F465",x"0E4A8",x"0DD0D",x"0D572",x"0C5B5",x"0C5D6",
									 x"0CE17",x"0CE79",x"0D6BA",x"0E73C",x"0F79E",x"0FFDF",x"0FFFF",x"1002A",x"0FFFF",x"1002D",
									 x"0F7BE",x"0EF5D",x"0E71B",x"0D69A",x"0C618",x"0BDF6",x"0C5D5",x"0D5B2",x"0D56F",x"0DCEA",
									 x"0E486",x"0EC84",x"0F4A3",x"0F4C3",x"0F4E2",x"0F503",x"0F524",x"0F544",x"0FD64",x"0FD84",
									 x"0FDA4",x"0FDC4",x"10000",x"0FDE4",x"10000",x"0FE04",x"0FE24",x"0FE25",x"0FE45",x"0FE44",
									 x"0FE45",x"0FE65",x"10001",x"0FE85",x"10003",x"0FEA5",x"10004",x"0FEC5",x"10006",x"0FEE5",
									 x"0FEE6",x"0FEE5",x"0FF05",x"0FF25",x"0FF46",x"10000",x"0FF65",x"0FF66",x"10000",x"0FF86",
									 x"0FFA6",x"10000",x"0FFC6",x"0FFA6",x"10000",x"0FFC7",x"10000",x"0FFA7",x"0FF87",x"0FF67",
									 x"0F767",x"10000",x"0F747",x"10001",x"0EF26",x"10003",x"0F746",x"10001",x"0F766",x"0F786",
									 x"0FFA7",x"10000",x"0FFC7",x"10001",x"0FFC6",x"0FFA6",x"0FFA7",x"10000",x"0FF86",x"10001",
									 x"0FF66",x"0FF45",x"0FF25",x"10000",x"0FF05",x"0FF06",x"10000",x"0FEC5",x"10001",x"0FEC6",
									 x"10002",x"0FEC5",x"10000",x"0FEA5",x"10004",x"0FE85",x"10002",x"0FE65",x"10002",x"0FE45",
									 x"10001",x"0FE25",x"0FE24",x"0FE04",x"10000",x"0FDE4",x"10000",x"0FDC4",x"0FDA4",x"10000",
									 x"0FD84",x"10000",x"0F564",x"0F544",x"0F503",x"0F4E3",x"0F4A3",x"0F482",x"0EC82",x"0E4A6",
									 x"0DCCA",x"0D52D",x"0CDB1",x"0CDF5",x"0C5F7",x"0C617",x"0CE79",x"0DEFB",x"0E73C",x"0F79E",
									 x"0FFFF",x"1002C",x"0FFFF",x"1002D",x"0FFDF",x"0F7BF",x"0EF7E",x"0E71C",x"0D69A",x"0C659",
									 x"0C617",x"0C5F6",x"0CDB5",x"0D570",x"0DCEB",x"0E4A7",x"0EC85",x"0F482",x"0FCA2",x"0FCC2",
									 x"0F4E3",x"0F523",x"0FD44",x"0FD64",x"0F584",x"10000",x"0F5A4",x"0FDA4",x"0FDC4",x"0FDE4",
									 x"10000",x"0FE04",x"10000",x"0FE24",x"0FE25",x"0FE45",x"10001",x"0FE65",x"10001",x"0FE85",
									 x"10003",x"0FEA5",x"10001",x"0FEC5",x"10006",x"0FEE6",x"0FEC6",x"0FEC5",x"10000",x"0FEE5",
									 x"0FF06",x"10000",x"0FF26",x"10000",x"0FF46",x"10000",x"0FF66",x"10000",x"0FF85",x"0FF86",
									 x"0FFA6",x"10003",x"0FFC6",x"0FFC7",x"10000",x"0FFA7",x"0FFC7",x"10005",x"0FFC6",x"10003",
									 x"0FFA6",x"0FFA7",x"10000",x"0FFA6",x"0FF86",x"10000",x"0FF65",x"0FF45",x"10000",x"0FF46",
									 x"0FF26",x"10000",x"0FF06",x"0FEE6",x"10004",x"0FEC5",x"10000",x"0FEC6",x"10003",x"0FEC5",
									 x"0FEA5",x"10003",x"0FE85",x"10003",x"0FE65",x"0FE45",x"10003",x"0FE24",x"10001",x"0FE04",
									 x"0FDE4",x"10000",x"0FDC4",x"0FDA4",x"10000",x"0FD84",x"0FD64",x"10000",x"0F544",x"0F523",
									 x"0F502",x"0F4C2",x"0F4A2",x"0F463",x"0F484",x"0ECC6",x"0DCEA",x"0D570",x"0CDB3",x"0C5F5",
									 x"0C617",x"0C638",x"0CE9A",x"0DF1B",x"0EF7D",x"0F79E",x"0FFDF",x"0FFFF",x"1002C",x"0FFFF",
									 x"1002E",x"0FFDF",x"0F7BF",x"0EF7E",x"0E71C",x"0D6BB",x"0CE39",x"0C5F8",x"0C5D7",x"0CDB5",
									 x"0D571",x"0DD0C",x"0E4A8",x"0F465",x"0FC63",x"0FC82",x"0F4C3",x"0F4E3",x"0F503",x"0FD24",
									 x"0FD64",x"0FD84",x"10000",x"0FDA4",x"10000",x"0FDC4",x"0FDE4",x"10000",x"0FE05",x"10000",
									 x"0FE25",x"10000",x"0FE45",x"10001",x"0FE65",x"10003",x"0FE85",x"10000",x"0FEA5",x"10005",
									 x"0FEC5",x"10003",x"0FEC6",x"10000",x"0FEE6",x"0FEE5",x"10000",x"0FEE6",x"10000",x"0FEE5",
									 x"0FF05",x"10001",x"0FF25",x"0FF26",x"0FF46",x"10002",x"0FF66",x"10000",x"0FF86",x"10001",
									 x"0FF87",x"10000",x"0FF86",x"10009",x"0FF66",x"0FF46",x"10000",x"0FF26",x"10002",x"0FF05",
									 x"10002",x"0FEE6",x"10000",x"0FEC5",x"10001",x"0FEC6",x"10002",x"0FEC5",x"0FEC6",x"10000",
									 x"0FEA6",x"10001",x"0FEA5",x"10000",x"0FE85",x"10003",x"0FE65",x"10000",x"0FE85",x"0FE65",
									 x"10000",x"0FE45",x"10000",x"0FE25",x"10002",x"0FE04",x"10000",x"0FDE4",x"0FDC4",x"10000",
									 x"0FDA4",x"10000",x"0F584",x"0FD64",x"0FD44",x"0FD24",x"0FD03",x"0FCE3",x"0FCC2",x"0FCA2",
									 x"0F483",x"0EC65",x"0EC87",x"0DCEB",x"0DD50",x"0CDB5",x"0C5F7",x"0BDF7",x"0CE59",x"0D6BA",
									 x"0DF1C",x"0EF7E",x"0F7DF",x"0FFDF",x"0FFFF",x"1002D",x"0FFFF",x"1002F",x"0FFDF",x"0F7BE",
									 x"0EF7D",x"0DF1C",x"0D6BA",x"0CE39",x"0BDF8",x"0C5D7",x"0CDB4",x"0CD92",x"0D52E",x"0DCCA",
									 x"0EC86",x"0EC64",x"0F483",x"0F4A3",x"0FCE3",x"0FD04",x"0FD24",x"0FD44",x"10000",x"0FD84",
									 x"10000",x"0FDA4",x"10000",x"0FDC4",x"0FDE4",x"0FE04",x"10001",x"0FE25",x"10000",x"0FE45",
									 x"10003",x"0FE65",x"10000",x"0FE85",x"10003",x"0FEA5",x"10002",x"0FEC5",x"10004",x"0FEE5",
									 x"10008",x"0FEE6",x"0FF06",x"10000",x"0FF26",x"10002",x"0FF46",x"1000B",x"0FF26",x"10004",
									 x"0FF06",x"10003",x"0FF05",x"0FF06",x"0FEE6",x"10000",x"0FEC5",x"10009",x"0FEA5",x"10001",
									 x"0FEA6",x"0FEA5",x"0FE85",x"10003",x"0FE65",x"10001",x"0FE45",x"10001",x"0FE25",x"10001",
									 x"0FE05",x"0FE04",x"10000",x"0FDE4",x"0FDC4",x"0FDA4",x"10001",x"0FD84",x"0FD64",x"0FD44",
									 x"0FD24",x"0FD04",x"0FCC3",x"0FCA3",x"0F483",x"0EC84",x"0E486",x"0DCCA",x"0DD0D",x"0CD71",
									 x"0CDB5",x"0C5D7",x"0C5F7",x"0C638",x"0D69A",x"0DEFC",x"0EF5D",x"0F7BE",x"0FFDF",x"0FFFF",
									 x"1002E",x"0FFFF",x"10031",x"0FFDF",x"0EFBE",x"0E75C",x"0DEDA",x"0CE9A",x"0C638",x"0C5F6",
									 x"0C5D5",x"0CDB4",x"0D550",x"0DCEC",x"0E4C8",x"0EC85",x"0F484",x"0FCA3",x"0FCC3",x"0FCE3",
									 x"0FD03",x"0FD23",x"0FD43",x"0FD63",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"0FDE4",x"10001",
									 x"0FE04",x"10000",x"0FE24",x"0FE25",x"0FE45",x"10002",x"0FE65",x"10000",x"0FE85",x"10002",
									 x"0FEA5",x"10005",x"0FEC5",x"10003",x"0FEE5",x"10000",x"0FEC5",x"10002",x"0FEE5",x"10003",
									 x"0FF05",x"10014",x"0FEE5",x"10004",x"0FEE6",x"10001",x"0FEC5",x"10009",x"0FEA5",x"10003",
									 x"0FE85",x"10003",x"0FE65",x"10000",x"0FE45",x"10001",x"0FE25",x"10001",x"0FE05",x"10000",
									 x"0FDE4",x"10000",x"0FDC4",x"10000",x"0FDA4",x"0FD84",x"10000",x"0FD63",x"0FD43",x"0FD23",
									 x"0F503",x"0FCE3",x"0F4C3",x"0F483",x"0F484",x"0EC85",x"0E4C8",x"0DCEB",x"0D52F",x"0CD92",
									 x"0C5F5",x"0C5F7",x"0CE39",x"0CE79",x"0D6BA",x"0E73C",x"0F77E",x"0FFBE",x"0FFFF",x"10030",
									 x"0FFFF",x"10033",x"0F7BE",x"0EF5C",x"0DEFB",x"0D6BA",x"0CE59",x"0BDF7",x"0C5D7",x"0CDD6",
									 x"0D593",x"0E52E",x"0E4CA",x"0EC67",x"0F464",x"0F482",x"10000",x"0FCC3",x"0F4E3",x"0FD03",
									 x"0FD24",x"0FD44",x"0FD64",x"0FD84",x"0FDA4",x"0FDC4",x"10000",x"0FDE4",x"10000",x"0FE04",
									 x"0FE05",x"10001",x"0FE25",x"10000",x"0FE45",x"10001",x"0FE65",x"10000",x"0FE85",x"10004",
									 x"0FEA5",x"10004",x"0FEC5",x"10004",x"0FEE5",x"10021",x"0FEC5",x"10004",x"0FEA5",x"10009",
									 x"0FE85",x"10003",x"0FE65",x"10000",x"0FE45",x"0FE44",x"10000",x"0FE24",x"10001",x"0FE05",
									 x"0FE04",x"0FDE5",x"10001",x"0FDC4",x"10000",x"0FDA4",x"0FD84",x"0FD64",x"0FD43",x"10000",
									 x"0FD03",x"0F4E3",x"10000",x"0F4C2",x"0F482",x"0F483",x"0ECA5",x"0E4C9",x"0DD2E",x"0D592",
									 x"0CDD5",x"0C5F6",x"0BDF7",x"0C638",x"0D6BA",x"0DEFB",x"0E73C",x"0F7BE",x"0FFFF",x"10032",
									 x"0FFFF",x"10034",x"0F79E",x"0EF5D",x"0E71C",x"0D6BA",x"0C658",x"0BDF7",x"10000",x"0C5D5",
									 x"0CD92",x"0D54F",x"0DCEA",x"0E4A6",x"0EC84",x"0F463",x"0F483",x"0F4C3",x"10000",x"0FCE4",
									 x"0FD04",x"0FD24",x"0FD44",x"0FD64",x"0FDA4",x"10000",x"0FDC4",x"10000",x"0FDE4",x"10001",
									 x"0FE05",x"10000",x"0FE25",x"10000",x"0FE45",x"10001",x"0FE65",x"10000",x"0FE85",x"10005",
									 x"0FEA5",x"10004",x"0FEC5",x"10003",x"0FEE5",x"1001A",x"0FEC5",x"1000A",x"0FEA5",x"10009",
									 x"0FE85",x"0FE65",x"10003",x"0FE45",x"10000",x"0FE24",x"10000",x"0FE04",x"10001",x"0FDE4",
									 x"10000",x"0FDC4",x"10001",x"0FDA4",x"10000",x"0FD84",x"0FD64",x"0FD23",x"10000",x"0F503",
									 x"0F4E4",x"0F4A3",x"0F483",x"0F482",x"0F484",x"0EC87",x"0DCCA",x"0D52D",x"0CD91",x"0C5B4",
									 x"0C5D6",x"0C5F7",x"0C618",x"0D69A",x"0DEFB",x"0E73C",x"0F79E",x"0FFDF",x"0FFFF",x"10032",
									 x"0FFFF",x"10034",x"0FFDF",x"0F7BE",x"0EF7D",x"0E73C",x"0D6DA",x"0CE79",x"0C638",x"0BDF7",
									 x"0C5F6",x"0CDD5",x"0CD91",x"0D50D",x"0E4A9",x"0EC87",x"0F465",x"0F4A3",x"10000",x"0FCC3",
									 x"0FCE3",x"0FD03",x"0FD23",x"0FD64",x"10000",x"0FD84",x"10000",x"0FDA4",x"0FDC4",x"10000",
									 x"0FDE4",x"10000",x"0FDE5",x"0FE05",x"0FE25",x"10001",x"0FE45",x"10000",x"0FE65",x"10001",
									 x"0FE85",x"10005",x"0FEA5",x"10003",x"0FEC5",x"10000",x"0FEA5",x"0FEC5",x"10008",x"0FEE5",
									 x"10010",x"0FEC5",x"1000A",x"0FEA5",x"10003",x"0FE85",x"10006",x"0FE65",x"10001",x"0FE45",
									 x"10001",x"0FE25",x"0FE24",x"0FE04",x"10001",x"0FDE4",x"0FDC4",x"10001",x"0FDA4",x"10000",
									 x"0FD84",x"0FD64",x"10000",x"0FD44",x"0FD03",x"0FCE3",x"10000",x"0F4C4",x"0F484",x"0F464",
									 x"0EC65",x"0E4A9",x"0DCED",x"0D551",x"0CDB3",x"0C5F5",x"0BDF6",x"0C617",x"0CE59",x"0D6BA",
									 x"0E71C",x"0EF7D",x"0F7BE",x"0FFDF",x"0FFFF",x"10033",x"0FFFF",x"10037",x"0F79E",x"0EF3C",
									 x"0E6FB",x"0D69B",x"0CE59",x"0C5F8",x"0C5D7",x"0C5B7",x"0CD95",x"0DD51",x"0E4ED",x"0E4A9",
									 x"0ECA6",x"0ECA4",x"0F483",x"0F4A2",x"0FCC2",x"0FCE2",x"0F503",x"0FD24",x"0FD44",x"0FD64",
									 x"0FD84",x"10000",x"0FDA4",x"10000",x"0FDC4",x"10000",x"0FDE4",x"10000",x"0FE04",x"10000",
									 x"0FE24",x"0FE25",x"0FE45",x"10000",x"0FE65",x"10002",x"0FE85",x"10000",x"0FE65",x"0FE85",
									 x"10001",x"0FEA5",x"10007",x"0FEC5",x"0FEA5",x"10000",x"0FEC5",x"10019",x"0FEA5",x"10007",
									 x"0FE85",x"10004",x"0FE65",x"10002",x"0FE45",x"10002",x"0FE24",x"10001",x"0FE05",x"0FE04",
									 x"0FDE4",x"10001",x"0FDC4",x"10000",x"0FDA4",x"0FD84",x"10000",x"0FD64",x"0FD44",x"0FD24",
									 x"0F503",x"0F4E3",x"0F4C3",x"0F4A3",x"10000",x"0F484",x"0F486",x"0ECA8",x"0DD0C",x"0D550",
									 x"0CD95",x"0C5B6",x"0BDD6",x"0BE18",x"0C659",x"0D69A",x"0E6FC",x"0E73C",x"0F79E",x"0FFDF",
									 x"0FFFF",x"10035",x"0FFFF",x"10037",x"0F7BE",x"0F79E",x"0EF5D",x"0E6FB",x"0D69A",x"0CE59",
									 x"0C618",x"0BDD9",x"0C5D7",x"0CDD5",x"0D592",x"0DD0E",x"0E4CA",x"0ECA7",x"0EC85",x"0F483",
									 x"0FCA3",x"0F4A2",x"0F4E3",x"0FD04",x"0FD24",x"0FD44",x"0FD64",x"10000",x"0FD84",x"0FDA4",
									 x"10000",x"0FDC4",x"10000",x"0FDE4",x"10000",x"0FE04",x"10000",x"0FE24",x"0FE25",x"0FE45",
									 x"10002",x"0FE65",x"10000",x"0FE45",x"0FE65",x"10002",x"0FE85",x"10002",x"0FEA5",x"1000A",
									 x"0FEC5",x"10014",x"0FEA5",x"10006",x"0FE85",x"10002",x"0FE65",x"10005",x"0FE45",x"10001",
									 x"0FE25",x"0FE24",x"0FE04",x"10000",x"0FE05",x"10000",x"0FDE4",x"0FDC4",x"10000",x"0FDA4",
									 x"10001",x"0FD84",x"0FD64",x"10000",x"0FD23",x"10000",x"0FD03",x"0FCE3",x"0F4C3",x"0F4A3",
									 x"0F483",x"0EC64",x"0E4A6",x"0DCCA",x"0D50D",x"0CD71",x"0CDD5",x"0BDF7",x"10000",x"0BE18",
									 x"0CE59",x"0D69A",x"0DEFB",x"0EF5D",x"0EF7D",x"0F7BE",x"0FFFF",x"10036",x"0FFFF",x"10038",
									 x"0FFDF",x"0F7BE",x"0EF7D",x"0E71B",x"0DEDA",x"0D679",x"0C638",x"0BE17",x"0BDF5",x"0BDB4",
									 x"0CD72",x"0DD30",x"0E4EC",x"0E4A8",x"0EC86",x"0F485",x"0F463",x"0F484",x"0F4C4",x"0F4E3",
									 x"0FD03",x"0FD23",x"0FD43",x"10000",x"0FD63",x"0F584",x"0FD84",x"0FDA4",x"0FDC4",x"10000",
									 x"0FDE4",x"10000",x"0FE04",x"10001",x"0FE24",x"10003",x"0FE44",x"0FE45",x"0FE65",x"10001",
									 x"0FE85",x"10004",x"0FEA5",x"10008",x"0FEC5",x"10010",x"0FEA5",x"1000A",x"0FE85",x"10000",
									 x"0FE65",x"10003",x"0FE45",x"10003",x"0FE25",x"0FE24",x"0FE04",x"10000",x"0FDE4",x"10002",
									 x"0FDC4",x"0FDA4",x"10001",x"0FD84",x"0FD64",x"0FD63",x"0FD43",x"0FD23",x"0FCE3",x"0FCC3",
									 x"0FCC2",x"0F4C2",x"0F4A3",x"0EC84",x"0EC85",x"0E4C7",x"0DD2C",x"0D56F",x"0CD72",x"0C5D4",
									 x"0C5F6",x"0BE17",x"0BE58",x"0CE99",x"0DEBA",x"0E6FB",x"0EF7D",x"0F7BE",x"0FFDF",x"0FFFF",
									 x"10037",x"0FFFF",x"1003A",x"0FFDF",x"0F7BE",x"0EF7D",x"0E71C",x"0D6DB",x"0CE7A",x"0C639",
									 x"0C618",x"0BDF7",x"0BDD6",x"0CDB3",x"0D550",x"0D4EC",x"0DCC9",x"0ECA6",x"0EC85",x"0EC83",
									 x"0F4A2",x"0F4E2",x"0FCE3",x"0F503",x"0FD03",x"0FD23",x"0FD44",x"0FD64",x"10000",x"0FD84",
									 x"0FD83",x"0FDA3",x"0FDA4",x"0FDC4",x"0FDE4",x"0FDE5",x"10000",x"0FE05",x"0FE04",x"10000",
									 x"0FE24",x"10002",x"0FE44",x"0FE45",x"10001",x"0FE65",x"10003",x"0FE85",x"10007",x"0FEA5",
									 x"10012",x"0FE85",x"10008",x"0FE65",x"10000",x"0FE45",x"0FE44",x"10001",x"0FE45",x"10001",
									 x"0FE25",x"10000",x"0FE05",x"0FE04",x"0FDE4",x"10000",x"0FDC4",x"10000",x"0FDC3",x"0FDA4",
									 x"10000",x"0FD83",x"0FD63",x"10000",x"0F544",x"0FD44",x"0FD23",x"0FD03",x"0FCE3",x"0FCC3",
									 x"0FCA3",x"0F4A3",x"0F483",x"0F484",x"0ECA6",x"0E4E9",x"0D50C",x"0CD50",x"0CD94",x"0C5D5",
									 x"0BDF7",x"0BE18",x"0C659",x"0CE79",x"0D6BA",x"0E73C",x"0EF7D",x"0F79E",x"0FFDF",x"0FFFF",
									 x"10039",x"0FFFF",x"1003B",x"0FFDF",x"0F7BE",x"0EF7D",x"0E73D",x"0DEDB",x"0D69A",x"0CE79",
									 x"0BDF7",x"0BDD6",x"0C5F7",x"0CDD6",x"0CD93",x"0DD50",x"0E4EB",x"0EC88",x"0F465",x"0F463",
									 x"0F4A2",x"10000",x"0F4A3",x"0F4C3",x"0F4E3",x"0F503",x"0FD04",x"0FD24",x"0FD44",x"0FD64",
									 x"0FD84",x"10000",x"0FDA4",x"0F5C4",x"10000",x"0FDE4",x"10002",x"0FE04",x"10000",x"0FE24",
									 x"10004",x"0FE45",x"10002",x"0FE65",x"10003",x"0FE85",x"1001B",x"0FE65",x"10004",x"0FE45",
									 x"0FE44",x"0FE24",x"10005",x"0FE04",x"0FE05",x"0FDE4",x"10002",x"0FDC4",x"0FDA4",x"10000",
									 x"0FD84",x"10000",x"0FD63",x"0FD42",x"0FD23",x"10000",x"0FD03",x"10000",x"0FCE3",x"0F4C3",
									 x"0F4A4",x"0F484",x"10000",x"0EC84",x"0E4A7",x"0DCEB",x"0D54F",x"0D593",x"0CDB4",x"0C5B6",
									 x"0BDB6",x"0BDF8",x"0C659",x"0D6BA",x"0DEDB",x"0E71C",x"0EF7D",x"0F7BE",x"0FFDF",x"0FFFF",
									 x"1003A",x"0FFFF",x"1003C",x"0FFDF",x"10000",x"0F79E",x"0EF3D",x"0DEFB",x"0D6BA",x"0CE59",
									 x"0C638",x"0C618",x"0C5F8",x"0BDD7",x"0C595",x"0D551",x"0DD0E",x"0ECAB",x"0ECA7",x"0ECA4",
									 x"0EC83",x"0F483",x"10000",x"0F4C3",x"0F4E3",x"0FCE3",x"0FD04",x"0FD24",x"10000",x"0FD44",
									 x"0FD64",x"0F584",x"0FDA4",x"10000",x"0FDC4",x"10002",x"0FDE4",x"10000",x"0FE04",x"10001",
									 x"0FE24",x"0FE25",x"10002",x"0FE24",x"10000",x"0FE45",x"10003",x"0FE65",x"10004",x"0FE85",
									 x"10010",x"0FE65",x"10004",x"0FE45",x"10004",x"0FE25",x"0FE24",x"10000",x"0FE04",x"10002",
									 x"0FDE4",x"10001",x"0FDC4",x"10002",x"0FDA4",x"10000",x"0FD84",x"0F564",x"0FD43",x"0F523",
									 x"0F522",x"0FD02",x"0FCE3",x"0FCC3",x"0FCC2",x"0FCA3",x"0F484",x"0EC85",x"0EC86",x"0ECA7",
									 x"0E4CA",x"0D50D",x"0CD51",x"0C5B4",x"0C5B6",x"0C5F7",x"0CE18",x"0C618",x"0CE59",x"0D6BB",
									 x"0E71B",x"0EF5C",x"0EF7D",x"0FFDF",x"0FFFF",x"1003C",x"0FFFF",x"1003E",x"0FFDF",x"0F79E",
									 x"0EF7D",x"0EF5D",x"0DEFB",x"0D6BA",x"0D678",x"0C617",x"0BDF7",x"0BDD7",x"0C5D6",x"0CDB4",
									 x"0D572",x"0D52E",x"0D4EA",x"0DCC7",x"0EC85",x"0F464",x"0EC83",x"0ECA3",x"0F4A3",x"0FCC3",
									 x"0FCE3",x"0F4E3",x"0F503",x"0FD24",x"0FD44",x"0FD64",x"10000",x"0FD84",x"10000",x"0FDA4",
									 x"10001",x"0FDC4",x"0FDE4",x"10005",x"0FE04",x"0FE05",x"10000",x"0FE25",x"10002",x"0FE45",
									 x"1000A",x"0FE65",x"10005",x"0FE45",x"1000B",x"0FE25",x"10003",x"0FE05",x"10000",x"0FDE4",
									 x"10001",x"0FDC4",x"10001",x"0FDA4",x"10001",x"0FD84",x"0FD83",x"0FD84",x"0FD64",x"0FD44",
									 x"0F524",x"0F523",x"0F503",x"10000",x"0F4E3",x"0F4C3",x"0F4A3",x"0F483",x"10000",x"0F484",
									 x"0EC86",x"0E488",x"0E4CA",x"0E50E",x"0DD52",x"0CD94",x"0C5D7",x"0C618",x"0BDF6",x"0C617",
									 x"0CE5A",x"0D69B",x"0DEFC",x"0E73D",x"0F79E",x"0F7BE",x"0FFDF",x"0FFFF",x"1003D",x"0FFFF",
									 x"10041",x"0FFDF",x"0EF9E",x"0EF5D",x"0E71B",x"0DEBA",x"0CE79",x"0C658",x"0BE17",x"0B5F7",
									 x"0BDD6",x"0C5B4",x"0CDB2",x"0D56F",x"0DD0D",x"0DCC9",x"0E4A7",x"0E486",x"0EC85",x"0F484",
									 x"0F4A3",x"10000",x"0F4C3",x"0F4E3",x"0FD03",x"10000",x"0FD23",x"0F543",x"10001",x"0F563",
									 x"0F583",x"10000",x"0FDA4",x"10002",x"0FDC4",x"10002",x"0FDE4",x"10001",x"0FE05",x"10004",
									 x"0FE25",x"10001",x"0FE24",x"10006",x"0FE45",x"0FE25",x"10001",x"0FE24",x"10004",x"0FE25",
									 x"10001",x"0FE05",x"10001",x"0FE25",x"0FE05",x"10002",x"0FDE4",x"10001",x"0FDC4",x"10001",
									 x"0FDA4",x"10002",x"0FD84",x"10000",x"0FD64",x"0FD44",x"0FD23",x"10001",x"0FD03",x"0F4E3",
									 x"10000",x"0F4C3",x"10000",x"0F4A3",x"0ECA4",x"0EC85",x"10000",x"0E487",x"0E4C9",x"0DD0D",
									 x"0D550",x"0D592",x"0CD94",x"0BDB6",x"0BDB7",x"0BDF8",x"0C638",x"0CE78",x"0D6BA",x"0E71C",
									 x"0EF5D",x"0EF7D",x"0F7BE",x"0FFFF",x"10040",x"0FFFF",x"10042",x"0FFBF",x"0FFBE",x"0EF7E",
									 x"0E73D",x"0DEFB",x"0D699",x"0C658",x"0BE38",x"0B5F7",x"0BDF7",x"0C5F7",x"0C5B6",x"0CD74",
									 x"0CD51",x"0DD0D",x"0E4AA",x"0EC88",x"0F486",x"0F464",x"0F484",x"0F483",x"0F4A3",x"0FCA3",
									 x"0FCC3",x"0FCE3",x"0F503",x"0F523",x"0F543",x"10001",x"0F563",x"0FD83",x"0FD84",x"10001",
									 x"0FDA4",x"10002",x"0FDC4",x"10001",x"0FDE4",x"10003",x"0FE04",x"0FE05",x"10001",x"0FE04",
									 x"10007",x"0FE24",x"10002",x"0FE04",x"10004",x"0FE05",x"0FE04",x"10000",x"0FDE4",x"10000",
									 x"0FDE5",x"0FDE4",x"10001",x"0FDC4",x"10002",x"0FDA4",x"10001",x"0FD83",x"10000",x"0FD84",
									 x"0FD64",x"0FD63",x"0F543",x"0FD43",x"0FD24",x"0FD03",x"0FCE3",x"10000",x"0FCC3",x"0F4C2",
									 x"0F4A2",x"0F4A3",x"0EC83",x"0ECA4",x"0ECA6",x"0ECA7",x"0E4EA",x"0DD2D",x"0D56F",x"0CD92",
									 x"0C5B5",x"0C5D7",x"0BDF8",x"0B618",x"0BE38",x"0C659",x"0D69A",x"0DEDB",x"0E71C",x"0F79D",
									 x"0F7BE",x"0FFDE",x"0FFFF",x"10041",x"0FFFF",x"10043",x"0FFDF",x"0F7BE",x"0F79E",x"0EF5D",
									 x"0E71C",x"0DEDB",x"0CE79",x"0C638",x"0BDF8",x"0BDD7",x"0BDB6",x"0C5B6",x"10000",x"0CD94",
									 x"0D550",x"0D50D",x"0DCCA",x"0E4A8",x"0EC87",x"0EC65",x"0F464",x"0F483",x"0FC83",x"0FCA3",
									 x"0F4C3",x"0FCE3",x"0FD03",x"10001",x"0FD23",x"0FD24",x"0FD44",x"10002",x"0FD64",x"10000",
									 x"0FD84",x"0FDA4",x"10001",x"0FDC4",x"10005",x"0FDC5",x"10001",x"0FDE5",x"10003",x"0FE05",
									 x"10004",x"0FDE5",x"10006",x"0FDC4",x"10003",x"0FDA4",x"10003",x"0FD84",x"10001",x"0FD64",
									 x"10000",x"0FD44",x"0FD43",x"0FD23",x"10000",x"0FD03",x"10000",x"0FCE3",x"0F4E3",x"0F4C3",
									 x"10000",x"0F4A3",x"0F483",x"0F482",x"0F463",x"0F484",x"0EC86",x"0E4A9",x"0DCCB",x"0D50D",
									 x"0CD50",x"0C5B3",x"0C5D5",x"0BDD6",x"10001",x"0C617",x"0C638",x"0CE79",x"0DEDB",x"0E71C",
									 x"0EF5D",x"0EF7D",x"0F7BE",x"0FFFF",x"10043",x"0FFFF",x"10045",x"0FFDF",x"0F7BE",x"0F79E",
									 x"0EF5D",x"0E71C",x"0D6DB",x"0CE79",x"0C658",x"0C638",x"0C617",x"0BDD6",x"0BDB5",x"0BD94",
									 x"0C593",x"0CD71",x"0D54F",x"0D50D",x"0DCCA",x"0E4A8",x"0ECA7",x"0EC85",x"0F484",x"10000",
									 x"0F4A4",x"0F4A3",x"0F4C3",x"0FCC3",x"0FCE3",x"10000",x"0FD03",x"0F503",x"0F523",x"0FD24",
									 x"10000",x"0FD44",x"10000",x"0FD64",x"10001",x"0FD84",x"0FD83",x"0FD84",x"0FDA4",x"10003",
									 x"0FDC4",x"10007",x"0FDE4",x"10002",x"0FDC4",x"10006",x"0FDA4",x"10003",x"0FD84",x"10002",
									 x"0FD63",x"0FD64",x"0FD44",x"0F544",x"0FD43",x"10000",x"0F523",x"0F503",x"0FD03",x"10000",
									 x"0F4E3",x"0F4C2",x"0F4A2",x"10000",x"0F4A3",x"0F4A4",x"0EC84",x"0EC85",x"0EC86",x"0E4A8",
									 x"0E4EA",x"0DD0C",x"0D54F",x"0CD71",x"0CD92",x"0C594",x"0C5B5",x"0C5D7",x"0C5F8",x"0C618",
									 x"0CE39",x"0D679",x"0D6BA",x"0E71C",x"0EF5D",x"0F79E",x"0F7BE",x"0FFDF",x"0FFFF",x"10044",
									 x"0FFFF",x"10048",x"0FFDF",x"0F79E",x"0EF5D",x"0E73C",x"0DEFB",x"0D6BA",x"0CE79",x"0C638",
									 x"0BE17",x"0B5F7",x"0BDF7",x"0C5D6",x"0C5B5",x"0C5B3",x"0CD70",x"0D52E",x"0DD0C",x"0E4EA",
									 x"0E4C8",x"0ECA7",x"0F4A6",x"0F485",x"0F484",x"0F4A3",x"0F4A2",x"0FCA2",x"0F4C2",x"10000",
									 x"0F4E2",x"0F503",x"10001",x"0FD23",x"0F523",x"0FD23",x"10000",x"0F543",x"0FD43",x"10001",
									 x"0FD63",x"0FD84",x"0FD83",x"0F584",x"0F5A4",x"0FD84",x"0FDA4",x"1000B",x"0FD84",x"0FDA4",
									 x"10002",x"0F583",x"10000",x"0FD83",x"0FD84",x"10000",x"0FD64",x"10000",x"0FD44",x"10000",
									 x"0FD43",x"10000",x"0F523",x"10000",x"0F503",x"10000",x"0FCE3",x"0F4E2",x"0FCE2",x"0FCC2",
									 x"0FCC3",x"0F4A3",x"10000",x"0F483",x"10000",x"0F4A5",x"0ECA6",x"0E4A8",x"0DCCB",x"0DCED",
									 x"0DD2F",x"0D551",x"0CD92",x"0C5D4",x"0BDF6",x"0C5F7",x"10000",x"0BDF7",x"0C619",x"0CE5A",
									 x"0D69A",x"0DEDB",x"0E71C",x"0EF5D",x"0EF7D",x"0FFDF",x"0FFFF",x"10047",x"0FFFF",x"10049",
									 x"0FFDF",x"0F7BE",x"0EF9E",x"0E75C",x"0DF1B",x"0D6DA",x"0CE9A",x"0C679",x"0C638",x"0BDF8",
									 x"0BDD7",x"0BDB6",x"0BDD5",x"0C5D5",x"0CDB4",x"0D5B3",x"0D550",x"0DD2E",x"0DCEC",x"0E4CA",
									 x"0ECA8",x"0EC87",x"0EC85",x"0EC84",x"0F483",x"10000",x"0F4A2",x"10000",x"0F4A3",x"0F4C2",
									 x"0FCC3",x"0FCE3",x"10000",x"0FD03",x"10000",x"0FD23",x"10001",x"0FD24",x"10000",x"0FD44",
									 x"0FD43",x"0F563",x"10000",x"0FD63",x"0FD64",x"10004",x"0FD84",x"0FD63",x"0FD84",x"10001",
									 x"0FD63",x"10005",x"0FD64",x"0F563",x"0FD44",x"10001",x"0FD24",x"10000",x"0FD23",x"0FD24",
									 x"0FD04",x"0FD03",x"0FCE3",x"10000",x"0FCC3",x"0FCA2",x"0F4A3",x"0F4A2",x"0F483",x"10000",
									 x"0F484",x"0EC84",x"0EC85",x"10000",x"0E487",x"0E4C9",x"0DCEB",x"0D50E",x"0D551",x"0D593",
									 x"0CD73",x"0CD94",x"0BDB5",x"0B5D6",x"0B5F7",x"0BE18",x"0C618",x"0C679",x"0D69A",x"0DEDB",
									 x"0DEFB",x"0EF5C",x"0F79D",x"0F7BE",x"0FFDF",x"0FFFF",x"10048",x"0FFFF",x"1004C",x"0F7BE",
									 x"0F79E",x"0EF7D",x"0E73C",x"0DEFB",x"0D69A",x"0CE79",x"0C638",x"0C618",x"0C5F8",x"0BDF7",
									 x"0BDD7",x"0C5D6",x"0C5B5",x"0C593",x"0CD72",x"0D551",x"0D52F",x"0D50D",x"0DCEB",x"0DCC9",
									 x"0E4A8",x"0E487",x"0EC85",x"10000",x"0EC84",x"0F484",x"0F483",x"10000",x"0F4A3",x"0F4C3",
									 x"10002",x"0F4E3",x"0F4E4",x"10000",x"0F504",x"0F503",x"10000",x"0F523",x"0FD03",x"0FD23",
									 x"10004",x"0FD24",x"0FD44",x"10002",x"0FD23",x"10000",x"0F503",x"0FD23",x"10002",x"0FD03",
									 x"0FD04",x"0F504",x"0FCE4",x"10000",x"0F4E4",x"10000",x"0F4C3",x"10000",x"0FCC3",x"0FCA3",
									 x"0F483",x"0F4A3",x"0F483",x"0F484",x"0EC84",x"0EC85",x"0EC86",x"0E4A7",x"0E4A8",x"0DCCA",
									 x"0DCCB",x"0DD0C",x"0D52E",x"0CD50",x"0CD71",x"0C573",x"0C5B4",x"0C5D6",x"10000",x"0C5F7",
									 x"0BDF7",x"0C618",x"0C638",x"0CE79",x"0D69A",x"0DEDB",x"0E71C",x"0EF5C",x"0F77D",x"0F7BE",
									 x"0FFFE",x"0FFFF",x"1004A",x"0FFFF",x"1004E",x"0FFDF",x"0F7BE",x"0F77E",x"0EF5D",x"0E71C",
									 x"0DEFB",x"0D6BA",x"0CE7A",x"0C639",x"0C618",x"0BE18",x"0B5D7",x"0BDD7",x"0BDD6",x"0C5D6",
									 x"0C5D5",x"0CDB4",x"0CD92",x"0D570",x"0D50E",x"0DCEC",x"0E4CA",x"0E4A9",x"0E4A8",x"0ECA7",
									 x"0EC86",x"0F485",x"0F484",x"10001",x"0F483",x"0F4A3",x"10000",x"0F4A4",x"0F4C4",x"0F4C3",
									 x"10004",x"0FCC3",x"10001",x"0F4C3",x"0F4E3",x"1000A",x"0F4C3",x"10001",x"0F4A3",x"0F4A4",
									 x"10003",x"0F484",x"0FC84",x"10000",x"0F484",x"0EC85",x"0ECA6",x"0ECA7",x"0E4C8",x"0E4E9",
									 x"0E4EB",x"0DD0D",x"0DD2E",x"0D570",x"0CD72",x"0CD94",x"0C5D5",x"10001",x"0BDD6",x"10000",
									 x"0BDF7",x"0BE18",x"0BE59",x"0CE7A",x"0D69A",x"0DEDB",x"0E71C",x"0E75C",x"0EF7E",x"0F79E",
									 x"0FFDF",x"10000",x"0FFFF",x"1004C",x"0FFFF",x"1004F",x"0FFDF",x"0F7BF",x"0F79E",x"0EF7D",
									 x"0EF5D",x"0E73C",x"0DEFB",x"0DEBA",x"0D67A",x"0CE59",x"0C638",x"10000",x"0BE18",x"0BE17",
									 x"0BDF6",x"0BDD6",x"0BDB5",x"0BD94",x"0C593",x"10000",x"0D572",x"0D551",x"0D52F",x"0DD2D",
									 x"0E4EC",x"0E4CA",x"0E4C9",x"0ECA8",x"0ECA7",x"0EC86",x"0F485",x"10000",x"0ECA5",x"10001",
									 x"0F4A4",x"0F484",x"0F483",x"0F4A3",x"10012",x"0ECA3",x"0F4A4",x"10001",x"0F484",x"10000",
									 x"0F485",x"0EC86",x"10000",x"0ECA7",x"0E4A9",x"0E4CA",x"0E4EC",x"0DD0D",x"0D52F",x"0D550",
									 x"0CD72",x"10000",x"0C573",x"0C594",x"0BDB5",x"0BDB6",x"0BDF6",x"0BE17",x"10000",x"0C637",
									 x"0C658",x"0CE79",x"0CE99",x"0D6BA",x"0DEFB",x"0E73C",x"0EF5C",x"0F77D",x"0F79D",x"0F7BE",
									 x"0FFDF",x"0FFFF",x"1004E",x"0FFFF",x"10050",x"0FFDF",x"10001",x"0F7BE",x"0F79E",x"0EF7D",
									 x"0E73C",x"0E6FC",x"0DEDB",x"0D6BA",x"0CE79",x"0C638",x"0C618",x"0BDF8",x"0BDD7",x"10000",
									 x"0BDB6",x"10001",x"0C5D6",x"0CDD5",x"0CD93",x"0CD92",x"0D571",x"0D54F",x"0D52E",x"0D50D",
									 x"0D4EC",x"0DCEB",x"0DCCA",x"0E4C9",x"0E4C7",x"0ECC7",x"0ECA6",x"0EC86",x"0EC85",x"0EC84",
									 x"0F483",x"10000",x"0F463",x"10001",x"0F462",x"10002",x"0F482",x"10001",x"0F462",x"10000",
									 x"0F463",x"0F483",x"10001",x"0EC64",x"0EC84",x"0EC85",x"0EC86",x"10000",x"0ECA7",x"0E4A8",
									 x"0E4C9",x"0DCCA",x"0DCCB",x"0D4EC",x"0D50D",x"0D52E",x"0D54F",x"0CD51",x"0CD72",x"0CD94",
									 x"0C5B4",x"0C5D5",x"0C5D6",x"0BDD6",x"10000",x"0BDD7",x"0BDF7",x"10000",x"0C618",x"0C638",
									 x"0CE79",x"0D6BA",x"0DEDB",x"0DEFB",x"0E73C",x"0EF7D",x"0F79D",x"0F7BE",x"0FFDE",x"0FFFF",
									 x"10051",x"0FFFF",x"10055",x"0FFDF",x"0F7BE",x"0F79E",x"0EF7D",x"0EF5D",x"0E73C",x"0E6FB",
									 x"0DEDB",x"0D6BB",x"0CE7A",x"0CE59",x"0C639",x"0C5F8",x"0BDF8",x"0BDF7",x"0B5D7",x"0BDD6",
									 x"0BDB5",x"10000",x"0BD94",x"0C594",x"0C593",x"0CD72",x"0CD71",x"0CD50",x"0D52E",x"0DD2C",
									 x"0DD0C",x"0E4EB",x"0E4CA",x"0E4C9",x"0E4A8",x"0E4A7",x"0E4A6",x"0E486",x"0EC86",x"0EC65",
									 x"10000",x"0EC64",x"10002",x"0EC84",x"0EC64",x"10000",x"0EC65",x"10000",x"0EC86",x"10000",
									 x"0E487",x"0E488",x"0E489",x"0E4A9",x"0E4CA",x"0DCCB",x"0DCEC",x"0DD0D",x"0D52E",x"0D550",
									 x"0CD71",x"0CD93",x"0C593",x"0BD94",x"10000",x"0BDB5",x"0BDB6",x"10000",x"0BDB7",x"0BDD7",
									 x"0BDF8",x"0BE18",x"0C639",x"0C659",x"0CE7A",x"0D69A",x"0DEDB",x"0E6DC",x"0E71C",x"0EF3D",
									 x"0EF5E",x"0F79E",x"0F7DF",x"10000",x"0FFFF",x"10054",x"0FFFF",x"10057",x"0F7DF",x"0F7DE",
									 x"0F7BE",x"0F77E",x"0EF5D",x"0EF3C",x"0E73C",x"0DEFB",x"0D6BA",x"0D69A",x"0CE79",x"0C659",
									 x"0C639",x"0BE18",x"10000",x"0C618",x"0BDF7",x"10001",x"0BDD6",x"0C5D5",x"0C5B4",x"0C593",
									 x"0C573",x"0C572",x"0C551",x"0CD30",x"0CD0F",x"10000",x"0CD0E",x"0CD0D",x"0D50D",x"10000",
									 x"0D4EC",x"10000",x"0D4EB",x"0D4CB",x"0DCEB",x"0DCEC",x"10002",x"0DCCB",x"10000",x"0D4CC",
									 x"0D4EC",x"0D4ED",x"10000",x"0CCEE",x"0CD0E",x"0CD0F",x"0CD2F",x"0CD30",x"0CD51",x"10000",
									 x"0CD72",x"0CD93",x"0C5B4",x"0C5D6",x"10000",x"0BDD7",x"10000",x"0BDF7",x"0BDF8",x"10000",
									 x"0C618",x"0C639",x"0C659",x"0CE79",x"0D69A",x"0DEBA",x"0DEDB",x"0E71C",x"0EF3D",x"0EF5D",
									 x"0F77E",x"0F79E",x"0FFBF",x"0FFDF",x"0FFFF",x"10056",x"0FFFF",x"1005A",x"0FFDF",x"0FFBF",
									 x"0F7BE",x"0F79D",x"0EF5D",x"0EF5C",x"0E73C",x"0DEFB",x"10000",x"0DEDA",x"0D69A",x"0CE79",
									 x"0CE59",x"0C658",x"0C638",x"0C618",x"0C617",x"0BDF7",x"0BDD6",x"0BDB5",x"0BD95",x"0B595",
									 x"10000",x"0BD95",x"0BD94",x"10000",x"0BD74",x"0BD93",x"0BD94",x"0C593",x"10000",x"0C573",
									 x"10002",x"0C593",x"10003",x"0C573",x"10000",x"0C574",x"10000",x"0C594",x"0BD94",x"0BD93",
									 x"0BD94",x"10001",x"0BD95",x"10000",x"0BDB5",x"0BDB6",x"0BDD6",x"0C5F7",x"0C617",x"0C618",
									 x"0C638",x"0CE58",x"0CE59",x"10000",x"0D699",x"0DEDA",x"0DEDB",x"0E6FB",x"0E71C",x"0EF3C",
									 x"0F75C",x"0F79D",x"0F79E",x"0F7BE",x"0FFDF",x"10000",x"0FFFF",x"10058",x"0FFFF",x"1005C",
									 x"0FFDF",x"10001",x"0FFBF",x"0F79E",x"0F77E",x"0F77D",x"0EF7D",x"0E73C",x"0E71C",x"10000",
									 x"0DEDB",x"0D6BA",x"10000",x"0CE99",x"0CE79",x"10000",x"0C659",x"0C639",x"0C618",x"0BE18",
									 x"0BDF7",x"10001",x"0BDD7",x"10005",x"0B5D7",x"10004",x"0BDD7",x"10003",x"0BDD8",x"0BDD7",
									 x"10000",x"0BDF7",x"0BDF8",x"10000",x"0BE18",x"0BE19",x"0C639",x"0C659",x"0CE59",x"0CE79",
									 x"0D699",x"0D69A",x"0D6BA",x"0DEDB",x"0DEFB",x"0E71C",x"0E73C",x"0EF5D",x"10000",x"0F79E",
									 x"0F7BE",x"0FFBF",x"0FFDF",x"0FFFF",x"1005D",x"0FFFF",x"10061",x"0FFDF",x"10001",x"0F79E",
									 x"10000",x"0EF7D",x"0EF5D",x"10000",x"0E73C",x"0E71C",x"0DEFB",x"10000",x"0DEDB",x"0D6BA",
									 x"10000",x"0CE79",x"0CE59",x"10000",x"0C638",x"10001",x"0C618",x"0BDF8",x"0BE18",x"0BDF8",
									 x"0BDF7",x"10005",x"0BDF8",x"10000",x"0C618",x"0BE18",x"0C618",x"10001",x"0C638",x"0C659",
									 x"0CE59",x"0CE79",x"0CE9A",x"0D69A",x"0D6BB",x"0DEDB",x"0DEFB",x"10000",x"0E71C",x"0E73C",
									 x"10000",x"0EF5D",x"0EF7D",x"0F79E",x"0F7BE",x"10000",x"0FFDF",x"0FFFF",x"10061",x"0FFFF",
									 x"10064",x"0FFDF",x"10001",x"0F7BE",x"0F79E",x"0EF7D",x"10001",x"0EF5D",x"0E73C",x"0E71C",
									 x"10000",x"0DEFB",x"0DEDB",x"10000",x"0D6BA",x"10000",x"0D69A",x"10000",x"0CE79",x"0D699",
									 x"0CE79",x"10003",x"0CE59",x"10000",x"0CE79",x"10003",x"0D69A",x"10001",x"0D6BA",x"10000",
									 x"0DEDB",x"10000",x"0DEFB",x"0E71C",x"10000",x"0E73C",x"0EF5D",x"10000",x"0EF7D",x"10000",
									 x"0F79E",x"0F7BE",x"0FFDF",x"10000",x"0FFFF",x"10064",x"0FFFF",x"10068",x"0FFDF",x"10001",
									 x"0F7BE",x"10000",x"0F79E",x"10000",x"0EF7D",x"10001",x"0EF5D",x"10000",x"0E73C",x"10000",
									 x"0E71C",x"10002",x"0DEFB",x"0E71C",x"0DEFB",x"10002",x"0E71C",x"0DEFB",x"10001",x"0E71C",
									 x"10001",x"0E73C",x"10000",x"0EF5D",x"10001",x"0EF7D",x"0F79E",x"10001",x"0F7BE",x"0FFDF",
									 x"10000",x"0FFFF",x"10069",x"0FFFF",x"1006F",x"0FFDF",x"10002",x"0F7BE",x"10000",x"0F79E",
									 x"10011",x"0F7BE",x"10000",x"0FFDF",x"10001",x"0FFFF",x"1006F",x"0FFFF",x"100FE",x"20008",
									 x"30000");

	------------------------------------------------------------------------------------------------
	-- Internal types	
	------------------------------------------------------------------------------------------------
	-- Define the different states of the statemachine	
	type compState is (normal, lineRepeatStart, lineRepeat, colRepeat, colLineRepeat);

	------------------------------------------------------------------------------------------------
	-- Internal signals	
	------------------------------------------------------------------------------------------------	
	-- Counter for the image signals
	signal cntH      : integer range 0 to imSizeH_g - 1;
	signal cntV      : integer range 0 to imSizeV_g - 1;
	
	-- Control signals for the image signals
	signal increment : std_logic;
	signal decrement : std_logic;

	-- Image signals
	signal color         : std_logic_vector(15 downto 0);
	signal valid        : std_logic;
	
	-- Signals for the deoding statemachine
	signal romCnt        : integer range 0 to (imSizeCompTotal_g);
	signal cntLineRepeat : integer range 0 to imSizeH_g - 1;
	signal cntColRepeat  : integer range 0 to imSizeV_g - 1;	
	signal oldColor      : std_logic_vector(15 downto 0);
	signal romCntSave    : integer range 0 to (imSizeCompTotal_g);
	signal romCntSaveLoc : integer range 0 to (imSizeCompTotal_g);
	signal curCompState : compState;

	-- ROM signals
	signal romData : std_logic_vector(17 downto 0);

begin
	-- Strobe out is set to the valid signal, which is set in the decoding statemachine
	strobe_out <= valid when resetn = '1' else '0';

	-- Set the image output signals
	row_out <= to_unsigned(cntH, rowSize_g);
	col_out <= to_unsigned(cntV, colSize_g);
	d_out   <= color;

	------------------------------------------------------------------------------------------------
	-- Read process
	------------------------------------------------------------------------------------------------
	rom_read : process(clk)
	begin
		-- Wait till the next rising edge occures
		if (rising_edge(clk)) then
			-- Read the requested data
			romData <= blockrom(romCnt);
		end if;
	end process rom_read;

	------------------------------------------------------------------------------------------------
	-- Row and Column process
	-- This process creates the signals to loop through all pixels
	------------------------------------------------------------------------------------------------
	changeRowColumn : process(clk)
	begin
		if rising_edge(clk) then
			if (resetn = '0') then
				-- Reset everything
				cntH       <= imSizeH_g - 1;
				cntV       <= imSizeV_g - 1;
				romCntSave <= 0;
			else
				-- Increment the row and column		
				if (increment = '1') then
					if (cntV = imSizeV_g - 1) then
						cntV <= 0;						
						if (cntH = imSizeH_g - 1) then
							cntH <= 0;
						else
							cntH <= cntH + 1;
						end if;
						
						-- We are on a new line - Save the current ROM address for the decoding statemachine
						if (romCnt > 0) then
							romCntSave <= romCnt - 1;
						else
							romCntSave <= 0;
						end if;
					else
						cntV <= cntV + 1;
					end if;
					
				-- Decrement the row and column					
				elsif (decrement = '1') then
					if (cntV = 0) then
						cntV <= imSizeV_g - 1;
						if (cntH = 0) then
							cntH <= imSizeH_g - 1;
						else
							cntH <= cntH - 1;
						end if;
					else
						cntV <= cntV - 1;
					end if;
				end if;
			end if;
		end if;
	end process changeRowColumn;

	------------------------------------------------------------------------------------------------
	-- Control process
	-- This process decodes the image
	------------------------------------------------------------------------------------------------
	control : process(clk)
	begin
		if rising_edge(clk) then
			if (resetn = '0') then
				-- Reset everything
				romCnt        <= 0;
				curCompState  <= normal;
				increment     <= '0';
				oldColor      <= (others => '0');
				cntColRepeat  <= 0;
				cntLineRepeat <= 0;
				romCntSaveLoc <= 0;
				decrement     <= '0';
				valid        <= '0';
			else
				-- Default assignements
				decrement <= '0';
				increment    <= '0';
				valid        <= '0';
				romCnt <= romCnt;
				curCompState <= curCompState;
				oldColor <= oldColor;
				cntColRepeat <= cntColRepeat;
				cntLineRepeat <= cntLineRepeat;
				romCntSaveLoc <= romCntSaveLoc;
				
				-- Statemachine
				case curCompState is
					-- No special decoding at the moment
					when normal =>						
						-- Decode command
						case romData(17 downto 16) is
							-- Repeat color command
							when "01" =>								
								cntColRepeat <= to_integer(unsigned(romData(15 downto 0)));
								curCompState <= colRepeat;								

							-- Repeat line command
							when "10" =>
								cntLineRepeat <= to_integer(unsigned(romData(15 downto 0)));
								romCntSaveLoc <= romCntSave;
								curCompState  <= lineRepeatStart;
								
							-- Normal color command
							when others =>
								increment <= '1';
								valid     <= '1';
								color     <= romData(15 downto 0);
								oldColor  <= romData(15 downto 0);
								
								if (romCnt = imSizeCompTotal_g - 1) then
									romCnt <= 0;
								else
									romCnt <= romCnt + 1;
								end if;
								
						end case;

					-- Execute color repeat command
					when colRepeat =>
						increment <= '1';
						valid     <= '1';
						color     <= oldColor;						
						
						if (cntColRepeat > 0) then
							cntColRepeat <= cntColRepeat - 1;
						else
							if (romCnt = imSizeCompTotal_g - 1) then
								romCnt <= 0;
							else
								romCnt <= romCnt + 1;
							end if;
							curCompState <= normal;
						end if;

					-- Execute line repeat command --> Is called at the start of a new line
					when lineRepeatStart =>
						decrement     <= '1';					
						cntLineRepeat <= cntLineRepeat - 1;
						romCnt        <= romCntSaveLoc;
						curCompState  <= lineRepeat;						

					-- Execute line repeat command 
					when lineRepeat =>
						if (cntV = imSizeV_g - 1) and (romCnt /= romCntSaveLoc + 1) then
							if (cntLineRepeat = 0) then
								curCompState <= normal;
								if (romCnt = imSizeCompTotal_g - 1) then
									romCnt <= 0;
								else
									romCnt <= romCnt + 1;
								end if;

							else
								curCompState <= lineRepeatStart;
							end if;

						else
							-- Decode command
							case romData(17 downto 16) is
								-- Repeat color command
								when "01" =>
									cntColRepeat <= to_integer(unsigned(romData(15 downto 0)));
									curCompState <= colLineRepeat;									

								-- Normal color command
								when others =>
									increment <= '1';
									valid     <= '1';
									color     <= romData(15 downto 0);
									oldColor  <= romData(15 downto 0);
									
									if (romCnt = imSizeCompTotal_g - 1) then
										romCnt <= 0;
									else
										romCnt <= romCnt + 1;
									end if;									
							end case;
						end if;

					-- Execute color repeat command during line repeat command
					when colLineRepeat =>						
						increment <= '1';
						valid     <= '1';
						color     <= oldColor;						
						
						if (cntColRepeat > 0) then
							cntColRepeat <= cntColRepeat - 1;
						else
							if (romCnt = imSizeCompTotal_g - 1) then
								romCnt <= 0;
							else
								romCnt <= romCnt + 1;
							end if;
							curCompState <= lineRepeat;
						end if;
				end case;
			end if;
		end if;
	end process control;
end architecture RTL;
